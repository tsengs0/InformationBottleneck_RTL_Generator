//`define SYM_CN_REV_1
//`define SYM_VN_REV_1
`define SYM_NO_IO_CONV
`define SHARED_ZERO_BS