module cnu6_ib_ram_wrapper #(
	parameter CN_ROM_RD_BW = 6,
	parameter CN_ROM_ADDR_BW = 10,
	parameter CN_PAGE_ADDR_BW = 5,
	parameter CN_DEGREE = 6,
	parameter IB_CNU_DECOMP_funNum = 4,
	parameter CN_NUM = 102,
	parameter CNU6_INSTANTIATE_NUM = 51,
	parameter CNU6_INSTANTIATE_UNIT = 2,
	parameter QUAN_SIZE = 4,
	parameter DATAPATH_WIDTH = 4
) (
	output wire read_addr_offset_out,
	output wire [DATAPATH_WIDTH-1:0] c2v_0_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_0_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_0_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_0_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_0_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_0_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_1_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_1_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_1_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_1_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_1_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_1_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_2_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_2_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_2_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_2_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_2_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_2_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_3_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_3_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_3_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_3_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_3_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_3_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_4_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_4_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_4_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_4_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_4_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_4_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_5_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_5_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_5_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_5_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_5_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_5_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_6_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_6_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_6_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_6_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_6_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_6_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_7_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_7_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_7_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_7_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_7_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_7_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_8_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_8_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_8_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_8_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_8_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_8_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_9_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_9_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_9_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_9_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_9_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_9_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_10_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_10_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_10_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_10_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_10_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_10_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_11_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_11_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_11_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_11_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_11_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_11_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_12_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_12_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_12_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_12_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_12_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_12_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_13_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_13_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_13_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_13_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_13_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_13_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_14_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_14_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_14_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_14_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_14_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_14_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_15_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_15_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_15_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_15_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_15_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_15_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_16_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_16_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_16_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_16_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_16_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_16_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_17_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_17_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_17_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_17_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_17_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_17_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_18_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_18_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_18_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_18_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_18_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_18_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_19_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_19_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_19_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_19_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_19_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_19_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_20_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_20_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_20_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_20_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_20_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_20_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_21_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_21_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_21_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_21_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_21_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_21_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_22_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_22_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_22_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_22_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_22_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_22_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_23_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_23_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_23_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_23_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_23_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_23_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_24_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_24_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_24_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_24_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_24_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_24_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_25_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_25_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_25_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_25_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_25_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_25_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_26_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_26_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_26_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_26_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_26_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_26_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_27_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_27_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_27_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_27_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_27_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_27_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_28_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_28_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_28_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_28_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_28_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_28_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_29_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_29_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_29_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_29_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_29_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_29_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_30_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_30_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_30_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_30_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_30_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_30_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_31_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_31_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_31_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_31_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_31_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_31_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_32_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_32_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_32_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_32_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_32_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_32_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_33_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_33_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_33_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_33_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_33_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_33_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_34_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_34_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_34_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_34_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_34_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_34_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_35_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_35_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_35_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_35_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_35_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_35_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_36_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_36_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_36_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_36_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_36_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_36_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_37_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_37_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_37_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_37_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_37_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_37_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_38_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_38_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_38_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_38_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_38_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_38_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_39_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_39_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_39_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_39_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_39_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_39_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_40_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_40_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_40_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_40_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_40_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_40_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_41_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_41_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_41_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_41_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_41_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_41_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_42_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_42_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_42_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_42_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_42_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_42_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_43_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_43_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_43_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_43_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_43_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_43_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_44_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_44_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_44_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_44_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_44_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_44_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_45_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_45_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_45_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_45_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_45_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_45_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_46_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_46_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_46_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_46_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_46_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_46_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_47_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_47_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_47_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_47_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_47_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_47_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_48_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_48_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_48_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_48_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_48_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_48_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_49_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_49_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_49_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_49_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_49_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_49_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_50_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_50_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_50_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_50_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_50_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_50_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_51_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_51_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_51_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_51_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_51_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_51_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_52_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_52_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_52_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_52_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_52_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_52_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_53_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_53_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_53_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_53_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_53_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_53_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_54_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_54_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_54_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_54_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_54_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_54_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_55_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_55_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_55_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_55_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_55_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_55_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_56_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_56_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_56_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_56_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_56_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_56_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_57_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_57_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_57_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_57_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_57_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_57_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_58_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_58_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_58_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_58_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_58_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_58_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_59_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_59_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_59_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_59_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_59_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_59_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_60_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_60_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_60_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_60_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_60_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_60_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_61_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_61_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_61_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_61_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_61_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_61_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_62_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_62_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_62_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_62_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_62_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_62_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_63_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_63_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_63_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_63_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_63_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_63_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_64_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_64_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_64_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_64_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_64_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_64_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_65_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_65_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_65_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_65_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_65_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_65_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_66_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_66_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_66_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_66_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_66_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_66_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_67_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_67_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_67_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_67_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_67_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_67_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_68_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_68_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_68_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_68_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_68_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_68_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_69_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_69_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_69_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_69_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_69_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_69_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_70_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_70_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_70_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_70_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_70_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_70_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_71_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_71_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_71_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_71_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_71_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_71_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_72_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_72_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_72_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_72_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_72_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_72_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_73_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_73_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_73_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_73_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_73_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_73_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_74_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_74_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_74_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_74_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_74_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_74_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_75_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_75_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_75_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_75_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_75_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_75_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_76_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_76_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_76_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_76_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_76_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_76_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_77_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_77_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_77_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_77_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_77_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_77_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_78_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_78_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_78_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_78_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_78_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_78_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_79_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_79_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_79_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_79_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_79_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_79_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_80_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_80_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_80_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_80_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_80_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_80_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_81_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_81_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_81_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_81_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_81_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_81_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_82_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_82_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_82_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_82_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_82_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_82_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_83_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_83_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_83_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_83_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_83_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_83_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_84_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_84_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_84_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_84_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_84_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_84_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_85_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_85_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_85_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_85_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_85_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_85_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_86_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_86_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_86_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_86_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_86_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_86_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_87_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_87_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_87_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_87_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_87_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_87_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_88_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_88_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_88_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_88_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_88_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_88_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_89_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_89_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_89_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_89_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_89_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_89_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_90_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_90_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_90_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_90_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_90_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_90_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_91_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_91_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_91_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_91_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_91_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_91_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_92_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_92_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_92_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_92_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_92_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_92_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_93_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_93_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_93_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_93_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_93_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_93_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_94_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_94_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_94_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_94_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_94_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_94_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_95_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_95_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_95_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_95_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_95_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_95_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_96_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_96_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_96_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_96_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_96_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_96_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_97_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_97_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_97_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_97_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_97_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_97_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_98_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_98_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_98_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_98_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_98_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_98_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_99_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_99_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_99_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_99_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_99_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_99_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_100_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_100_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_100_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_100_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_100_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_100_out5,
	output wire [DATAPATH_WIDTH-1:0] c2v_101_out0,
	output wire [DATAPATH_WIDTH-1:0] c2v_101_out1,
	output wire [DATAPATH_WIDTH-1:0] c2v_101_out2,
	output wire [DATAPATH_WIDTH-1:0] c2v_101_out3,
	output wire [DATAPATH_WIDTH-1:0] c2v_101_out4,
	output wire [DATAPATH_WIDTH-1:0] c2v_101_out5,

	input wire [DATAPATH_WIDTH-1:0] v2c_0_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_0_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_0_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_0_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_0_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_0_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_1_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_1_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_1_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_1_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_1_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_1_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_2_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_2_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_2_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_2_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_2_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_2_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_3_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_3_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_3_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_3_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_3_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_3_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_4_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_4_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_4_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_4_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_4_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_4_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_5_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_5_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_5_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_5_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_5_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_5_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_6_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_6_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_6_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_6_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_6_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_6_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_7_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_7_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_7_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_7_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_7_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_7_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_8_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_8_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_8_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_8_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_8_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_8_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_9_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_9_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_9_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_9_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_9_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_9_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_10_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_10_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_10_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_10_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_10_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_10_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_11_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_11_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_11_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_11_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_11_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_11_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_12_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_12_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_12_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_12_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_12_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_12_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_13_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_13_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_13_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_13_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_13_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_13_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_14_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_14_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_14_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_14_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_14_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_14_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_15_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_15_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_15_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_15_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_15_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_15_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_16_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_16_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_16_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_16_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_16_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_16_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_17_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_17_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_17_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_17_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_17_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_17_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_18_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_18_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_18_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_18_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_18_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_18_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_19_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_19_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_19_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_19_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_19_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_19_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_20_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_20_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_20_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_20_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_20_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_20_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_21_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_21_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_21_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_21_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_21_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_21_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_22_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_22_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_22_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_22_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_22_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_22_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_23_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_23_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_23_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_23_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_23_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_23_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_24_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_24_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_24_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_24_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_24_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_24_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_25_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_25_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_25_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_25_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_25_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_25_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_26_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_26_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_26_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_26_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_26_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_26_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_27_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_27_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_27_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_27_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_27_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_27_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_28_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_28_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_28_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_28_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_28_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_28_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_29_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_29_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_29_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_29_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_29_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_29_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_30_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_30_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_30_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_30_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_30_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_30_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_31_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_31_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_31_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_31_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_31_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_31_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_32_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_32_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_32_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_32_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_32_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_32_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_33_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_33_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_33_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_33_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_33_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_33_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_34_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_34_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_34_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_34_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_34_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_34_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_35_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_35_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_35_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_35_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_35_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_35_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_36_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_36_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_36_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_36_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_36_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_36_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_37_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_37_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_37_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_37_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_37_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_37_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_38_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_38_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_38_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_38_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_38_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_38_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_39_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_39_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_39_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_39_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_39_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_39_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_40_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_40_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_40_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_40_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_40_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_40_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_41_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_41_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_41_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_41_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_41_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_41_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_42_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_42_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_42_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_42_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_42_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_42_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_43_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_43_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_43_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_43_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_43_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_43_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_44_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_44_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_44_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_44_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_44_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_44_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_45_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_45_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_45_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_45_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_45_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_45_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_46_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_46_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_46_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_46_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_46_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_46_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_47_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_47_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_47_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_47_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_47_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_47_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_48_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_48_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_48_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_48_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_48_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_48_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_49_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_49_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_49_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_49_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_49_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_49_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_50_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_50_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_50_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_50_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_50_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_50_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_51_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_51_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_51_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_51_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_51_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_51_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_52_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_52_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_52_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_52_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_52_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_52_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_53_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_53_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_53_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_53_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_53_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_53_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_54_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_54_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_54_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_54_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_54_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_54_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_55_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_55_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_55_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_55_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_55_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_55_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_56_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_56_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_56_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_56_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_56_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_56_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_57_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_57_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_57_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_57_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_57_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_57_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_58_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_58_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_58_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_58_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_58_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_58_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_59_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_59_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_59_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_59_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_59_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_59_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_60_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_60_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_60_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_60_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_60_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_60_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_61_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_61_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_61_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_61_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_61_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_61_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_62_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_62_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_62_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_62_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_62_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_62_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_63_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_63_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_63_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_63_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_63_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_63_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_64_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_64_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_64_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_64_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_64_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_64_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_65_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_65_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_65_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_65_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_65_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_65_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_66_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_66_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_66_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_66_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_66_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_66_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_67_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_67_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_67_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_67_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_67_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_67_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_68_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_68_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_68_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_68_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_68_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_68_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_69_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_69_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_69_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_69_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_69_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_69_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_70_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_70_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_70_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_70_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_70_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_70_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_71_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_71_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_71_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_71_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_71_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_71_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_72_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_72_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_72_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_72_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_72_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_72_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_73_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_73_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_73_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_73_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_73_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_73_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_74_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_74_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_74_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_74_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_74_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_74_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_75_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_75_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_75_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_75_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_75_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_75_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_76_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_76_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_76_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_76_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_76_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_76_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_77_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_77_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_77_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_77_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_77_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_77_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_78_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_78_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_78_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_78_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_78_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_78_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_79_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_79_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_79_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_79_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_79_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_79_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_80_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_80_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_80_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_80_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_80_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_80_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_81_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_81_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_81_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_81_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_81_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_81_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_82_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_82_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_82_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_82_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_82_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_82_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_83_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_83_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_83_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_83_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_83_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_83_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_84_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_84_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_84_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_84_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_84_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_84_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_85_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_85_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_85_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_85_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_85_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_85_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_86_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_86_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_86_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_86_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_86_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_86_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_87_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_87_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_87_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_87_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_87_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_87_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_88_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_88_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_88_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_88_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_88_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_88_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_89_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_89_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_89_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_89_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_89_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_89_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_90_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_90_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_90_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_90_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_90_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_90_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_91_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_91_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_91_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_91_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_91_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_91_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_92_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_92_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_92_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_92_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_92_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_92_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_93_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_93_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_93_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_93_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_93_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_93_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_94_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_94_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_94_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_94_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_94_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_94_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_95_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_95_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_95_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_95_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_95_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_95_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_96_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_96_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_96_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_96_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_96_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_96_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_97_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_97_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_97_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_97_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_97_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_97_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_98_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_98_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_98_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_98_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_98_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_98_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_99_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_99_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_99_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_99_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_99_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_99_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_100_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_100_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_100_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_100_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_100_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_100_in5,
	input wire [DATAPATH_WIDTH-1:0] v2c_101_in0,
	input wire [DATAPATH_WIDTH-1:0] v2c_101_in1,
	input wire [DATAPATH_WIDTH-1:0] v2c_101_in2,
	input wire [DATAPATH_WIDTH-1:0] v2c_101_in3,
	input wire [DATAPATH_WIDTH-1:0] v2c_101_in4,
	input wire [DATAPATH_WIDTH-1:0] v2c_101_in5,

	input wire read_clk,
	input wire read_addr_offset,
	input wire v2c_latch_en,
	input wire v2c_parallel_load,

	// Iteration-Refresh Page Address
	input wire [CN_PAGE_ADDR_BW+1-1:0] page_addr_ram_0,
	input wire [CN_PAGE_ADDR_BW+1-1:0] page_addr_ram_1,
	input wire [CN_PAGE_ADDR_BW+1-1:0] page_addr_ram_2,
	input wire [CN_PAGE_ADDR_BW+1-1:0] page_addr_ram_3,
	//Iteration-Refresh Page Data
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataA_0, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataB_0, // from portB of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataA_1, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataB_1, // from portB of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataA_2, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataB_2, // from portB of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataA_3, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] ram_write_dataB_3, // from portB of IB-ROM

	input wire [3:0] ib_ram_we,
	input wire write_clk
);
// Input sources of check node units
wire [QUAN_SIZE-1:0] v2c_0 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] v2c_1 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] v2c_2 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] v2c_3 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] v2c_4 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] v2c_5 [0:CN_NUM-1];
// Output sources of check node units
wire [QUAN_SIZE-1:0] c2v_0 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] c2v_1 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] c2v_2 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] c2v_3 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] c2v_4 [0:CN_NUM-1];
wire [QUAN_SIZE-1:0] c2v_5 [0:CN_NUM-1];
// Address related signals including the Net type
wire [CN_DEGREE-2-1-1:0] read_addr_offset_internal [0:CNU6_INSTANTIATE_NUM-1];
wire [CNU6_INSTANTIATE_NUM-1:0]read_addr_offset_outSet;

reg [DATAPATH_WIDTH-1:0] v2c_latch_0 [0:CN_NUM-1];
reg [DATAPATH_WIDTH-1:0] v2c_latch_1 [0:CN_NUM-1];
reg [DATAPATH_WIDTH-1:0] v2c_latch_2 [0:CN_NUM-1];
reg [DATAPATH_WIDTH-1:0] v2c_latch_3 [0:CN_NUM-1];
reg [DATAPATH_WIDTH-1:0] v2c_latch_4 [0:CN_NUM-1];
reg [DATAPATH_WIDTH-1:0] v2c_latch_5 [0:CN_NUM-1];
generate 
	genvar j;
	for (j=0; j<CNU6_INSTANTIATE_NUM; j=j+1) begin : v2c_latch_inst
	///////////////////////////////////////////////////////////////////////////////////////////
	// v2c_out_0
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_0[(CNU6_INSTANTIATE_UNIT*j)];
		else 
			v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)];
	end
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)+1] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_0[(CNU6_INSTANTIATE_UNIT*j)+1];
		else 
			v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)+1];
	end	
	///////////////////////////////////////////////////////////////////////////////////////////
	// v2c_out_1
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_1[(CNU6_INSTANTIATE_UNIT*j)];
		else 
			v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)];
	end
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)+1] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_1[(CNU6_INSTANTIATE_UNIT*j)+1];
		else 
			v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)+1];
	end	
	///////////////////////////////////////////////////////////////////////////////////////////
	// v2c_out_2
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_2[(CNU6_INSTANTIATE_UNIT*j)];
		else 
			v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)];
	end
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)+1] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_2[(CNU6_INSTANTIATE_UNIT*j)+1];
		else 
			v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)+1];
	end	
	///////////////////////////////////////////////////////////////////////////////////////////
	// v2c_out_3
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_3[(CNU6_INSTANTIATE_UNIT*j)];
		else 
			v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)];
	end
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)+1] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_3[(CNU6_INSTANTIATE_UNIT*j)+1];
		else 
			v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)+1];
	end	
	///////////////////////////////////////////////////////////////////////////////////////////
	// v2c_out_4
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_4[(CNU6_INSTANTIATE_UNIT*j)];
		else 
			v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)];
	end
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)+1] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_4[(CNU6_INSTANTIATE_UNIT*j)+1];
		else 
			v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)+1];
	end	
	///////////////////////////////////////////////////////////////////////////////////////////
	// v2c_out_5
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_5[(CNU6_INSTANTIATE_UNIT*j)];
		else 
			v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)] <= v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)];
	end
	always @(posedge read_clk, posedge v2c_latch_en) begin
		if(v2c_parallel_load == 1'b1) // from v2c_load[0]
			v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)+1] <= 0;
		else if(v2c_latch_en == 1'b1) 
			v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_5[(CNU6_INSTANTIATE_UNIT*j)+1];
		else 
			v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)+1] <= v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)+1];
	end	
	///////////////////////////////////////////////////////////////////////////////////////////
end
endgenerate

generate
  //genvar j;
  // Group A interacting with Port A of IB-ROMs
  localparam inst_num_groupA = 25;  
  for (j=0; j<inst_num_groupA; j=j+1) begin : cnu6_204_102_inst_GroupA
    // Instantiation of F_0
    wire [QUAN_SIZE-1:0] f0_out[0:3];
    wire [QUAN_SIZE-1:0] cnu0_f0_M_reg [0:CN_DEGREE-1];
    wire [QUAN_SIZE-1:0] cnu1_f0_M_reg [0:CN_DEGREE-1];
		
    cnu6_f0 u_f0(
		.read_addr_offset_out (read_addr_offset_internal[j][0]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .t_portA (f0_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portB (f0_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        // For the second CNU
        .t_portC (f0_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portD (f0_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the first CNU
        .cnu0_M_reg0 (cnu0_f0_M_reg[0]),
        .cnu0_M_reg1 (cnu0_f0_M_reg[1]),
        .cnu0_M_reg2 (cnu0_f0_M_reg[2]),
        .cnu0_M_reg3 (cnu0_f0_M_reg[3]),
        .cnu0_M_reg4 (cnu0_f0_M_reg[4]),
        .cnu0_M_reg5 (cnu0_f0_M_reg[5]),
        // For the second CNU
        .cnu1_M_reg0 (cnu1_f0_M_reg[0]),
        .cnu1_M_reg1 (cnu1_f0_M_reg[1]),
        .cnu1_M_reg2 (cnu1_f0_M_reg[2]),
        .cnu1_M_reg3 (cnu1_f0_M_reg[3]),
        .cnu1_M_reg4 (cnu1_f0_M_reg[4]),
        .cnu1_M_reg5 (cnu1_f0_M_reg[5]),

        // From the first CNU
        .cnu0_v2c_0 (/*v2c_0*/v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_1 (/*v2c_1*/v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_2 (/*v2c_2*/v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_3 (/*v2c_3*/v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_4 (/*v2c_4*/v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_5 (/*v2c_5*/v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)]),
        // From the second CNU
        .cnu1_v2c_0 (/*v2c_0*/v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_1 (/*v2c_1*/v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_2 (/*v2c_2*/v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_3 (/*v2c_3*/v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_4 (/*v2c_4*/v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_5 (/*v2c_5*/v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)+1]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset), // offset determing the switch between multi-frame under the following sub-datapath
	
		// Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_0[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_0 (ram_write_dataA_0[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[0])
    );
    // Instantiation of F_1
    wire [QUAN_SIZE-1:0] f1_out[0:3];
    wire [QUAN_SIZE-1:0] cnu0_f1_M_reg [0:CN_DEGREE-1];
    wire [QUAN_SIZE-1:0] cnu1_f1_M_reg [0:CN_DEGREE-1];
    cnu6_f1 u_f1(
		.read_addr_offset_out (read_addr_offset_internal[j][1]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .t_portA (f1_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portB (f1_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        // For the second CNU
        .t_portC (f1_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portD (f1_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the first CNU
        .cnu0_M_reg0 (cnu0_f1_M_reg[0]),
        .cnu0_M_reg1 (cnu0_f1_M_reg[1]),
        .cnu0_M_reg2 (cnu0_f1_M_reg[2]),
        .cnu0_M_reg3 (cnu0_f1_M_reg[3]),
        .cnu0_M_reg4 (cnu0_f1_M_reg[4]),
        .cnu0_M_reg5 (cnu0_f1_M_reg[5]),
        // For the second CNU
        .cnu1_M_reg0 (cnu1_f1_M_reg[0]),
        .cnu1_M_reg1 (cnu1_f1_M_reg[1]),
        .cnu1_M_reg2 (cnu1_f1_M_reg[2]),
        .cnu1_M_reg3 (cnu1_f1_M_reg[3]),
        .cnu1_M_reg4 (cnu1_f1_M_reg[4]),
        .cnu1_M_reg5 (cnu1_f1_M_reg[5]),

        // From the first CNU
        .t_00 (f0_out[0]),
        .t_01 (f0_out[1]),
        .cnu0_v2c_0 (cnu0_f0_M_reg[0]),
        .cnu0_v2c_1 (cnu0_f0_M_reg[1]),
        .cnu0_v2c_2 (cnu0_f0_M_reg[2]),
        .cnu0_v2c_3 (cnu0_f0_M_reg[3]),
        .cnu0_v2c_4 (cnu0_f0_M_reg[4]),
        .cnu0_v2c_5 (cnu0_f0_M_reg[5]),
        // From the second CNU
        .t_02 (f0_out[2]),
        .t_03 (f0_out[3]),
        .cnu1_v2c_0 (cnu1_f0_M_reg[0]),
        .cnu1_v2c_1 (cnu1_f0_M_reg[1]),
        .cnu1_v2c_2 (cnu1_f0_M_reg[2]),
        .cnu1_v2c_3 (cnu1_f0_M_reg[3]),
        .cnu1_v2c_4 (cnu1_f0_M_reg[4]),
        .cnu1_v2c_5 (cnu1_f0_M_reg[5]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset_internal[j][0]), // offset determing the switch between multi-frame under the following sub-datapath

        // Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_1[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_1 (ram_write_dataA_1[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[1])
    );
    // Instantiation of F_2
    wire [QUAN_SIZE-1:0] cnu0_f2_out[0:3];
    wire [QUAN_SIZE-1:0] cnu1_f2_out[0:3];
    wire [QUAN_SIZE-1:0] cnu0_f2_M_reg [0:3];
    wire [QUAN_SIZE-1:0] cnu1_f2_M_reg [0:3];
    cnu6_f2 u_f2(
		.read_addr_offset_out (read_addr_offset_internal[j][2]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .cnu0_t_portA (cnu0_f2_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu0_t_portB (cnu0_f2_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu0_t_portC (cnu0_f2_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu0_t_portD (cnu0_f2_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the second CNU
        .cnu1_t_portA (cnu1_f2_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu1_t_portB (cnu1_f2_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu1_t_portC (cnu1_f2_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu1_t_portD (cnu1_f2_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the first CNU
        .cnu0_M_reg1 (cnu0_f2_M_reg[0]),
        .cnu0_M_reg2 (cnu0_f2_M_reg[1]),
        .cnu0_M_reg4 (cnu0_f2_M_reg[2]),
        .cnu0_M_reg5 (cnu0_f2_M_reg[3]),
        // For the second CNU
        .cnu1_M_reg1 (cnu1_f2_M_reg[0]),
        .cnu1_M_reg2 (cnu1_f2_M_reg[1]),
        .cnu1_M_reg4 (cnu1_f2_M_reg[2]),
        .cnu1_M_reg5 (cnu1_f2_M_reg[3]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset_internal[j][1]), // offset determing the switch between multi-frame under the following sub-datapath

        // From the first CNU
        .t_10 (f1_out[0]),
        .t_11 (f1_out[1]),
        .cnu0_v2c_0 (cnu0_f1_M_reg[0]),
        .cnu0_v2c_1 (cnu0_f1_M_reg[1]),
        .cnu0_v2c_2 (cnu0_f1_M_reg[2]),
        .cnu0_v2c_3 (cnu0_f1_M_reg[3]),
        .cnu0_v2c_4 (cnu0_f1_M_reg[4]),
        .cnu0_v2c_5 (cnu0_f1_M_reg[5]),
        // From the second CNU
        .t_12 (f1_out[2]),
        .t_13 (f1_out[3]),
        .cnu1_v2c_0 (cnu1_f1_M_reg[0]),
        .cnu1_v2c_1 (cnu1_f1_M_reg[1]),
        .cnu1_v2c_2 (cnu1_f1_M_reg[2]),
        .cnu1_v2c_3 (cnu1_f1_M_reg[3]),
        .cnu1_v2c_4 (cnu1_f1_M_reg[4]),
        .cnu1_v2c_5 (cnu1_f1_M_reg[5]),

        // Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_2[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_2 (ram_write_dataA_2[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[2])
    );
    // Instantiation of F_3
    wire [QUAN_SIZE-1:0] cnu0_c2v [0:CN_DEGREE-1];
    wire [QUAN_SIZE-1:0] cnu1_c2v [0:CN_DEGREE-1];
    cnu6_f3 u_f3(
		.read_addr_offset_out (read_addr_offset_outSet[j]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .cnu0_c2v_0 (c2v_0[(CNU6_INSTANTIATE_UNIT*j)]), 
        .cnu0_c2v_1 (c2v_1[(CNU6_INSTANTIATE_UNIT*j)]), 
        .cnu0_c2v_2 (c2v_2[(CNU6_INSTANTIATE_UNIT*j)]), 
        .cnu0_c2v_3 (c2v_3[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_c2v_4 (c2v_4[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_c2v_5 (c2v_5[(CNU6_INSTANTIATE_UNIT*j)]), 
        // For the second CNU
        .cnu1_c2v_0 (c2v_0[(CNU6_INSTANTIATE_UNIT*j)+1]), 
        .cnu1_c2v_1 (c2v_1[(CNU6_INSTANTIATE_UNIT*j)+1]), 
        .cnu1_c2v_2 (c2v_2[(CNU6_INSTANTIATE_UNIT*j)+1]), 
        .cnu1_c2v_3 (c2v_3[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_c2v_4 (c2v_4[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_c2v_5 (c2v_5[(CNU6_INSTANTIATE_UNIT*j)+1]),

        // From the first CNU
        .cnu0_t_20 (cnu0_f2_out[0]),
        .cnu0_t_21 (cnu0_f2_out[1]),
        .cnu0_t_22 (cnu0_f2_out[2]),
        .cnu0_t_23 (cnu0_f2_out[3]),
        .cnu0_v2c_1 (cnu0_f2_M_reg[0]),
        .cnu0_v2c_2 (cnu0_f2_M_reg[1]),
        .cnu0_v2c_4 (cnu0_f2_M_reg[2]),
        .cnu0_v2c_5 (cnu0_f2_M_reg[3]),
        // From the second CNU
        .cnu1_t_20 (cnu1_f2_out[0]),
        .cnu1_t_21 (cnu1_f2_out[1]),
        .cnu1_t_22 (cnu1_f2_out[2]),
        .cnu1_t_23 (cnu1_f2_out[3]),
        .cnu1_v2c_1 (cnu1_f2_M_reg[0]),
        .cnu1_v2c_2 (cnu1_f2_M_reg[1]),
        .cnu1_v2c_4 (cnu1_f2_M_reg[2]),
        .cnu1_v2c_5 (cnu1_f2_M_reg[3]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset_internal[j][2]), // offset determing the switch between multi-frame under the following sub-datapath

        // Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_3[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_3 (ram_write_dataA_3[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[3])
    );
  end
  
   // Group B interacting with Port B of IB-ROMs
   localparam inst_num_groupB = 26;
   for (j=inst_num_groupB-1; j<CNU6_INSTANTIATE_NUM; j=j+1) begin : cnu6_204_102_inst_GroupB
    // Instantiation of F_0
    wire [QUAN_SIZE-1:0] f0_out[0:3];
    wire [QUAN_SIZE-1:0] cnu0_f0_M_reg [0:CN_DEGREE-1];
    wire [QUAN_SIZE-1:0] cnu1_f0_M_reg [0:CN_DEGREE-1];
    cnu6_f0 u_f0(
		.read_addr_offset_out (read_addr_offset_internal[j][0]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .t_portA (f0_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portB (f0_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        // For the second CNU
        .t_portC (f0_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portD (f0_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the first CNU
        .cnu0_M_reg0 (cnu0_f0_M_reg[0]),
        .cnu0_M_reg1 (cnu0_f0_M_reg[1]),
        .cnu0_M_reg2 (cnu0_f0_M_reg[2]),
        .cnu0_M_reg3 (cnu0_f0_M_reg[3]),
        .cnu0_M_reg4 (cnu0_f0_M_reg[4]),
        .cnu0_M_reg5 (cnu0_f0_M_reg[5]),
        // For the second CNU
        .cnu1_M_reg0 (cnu1_f0_M_reg[0]),
        .cnu1_M_reg1 (cnu1_f0_M_reg[1]),
        .cnu1_M_reg2 (cnu1_f0_M_reg[2]),
        .cnu1_M_reg3 (cnu1_f0_M_reg[3]),
        .cnu1_M_reg4 (cnu1_f0_M_reg[4]),
        .cnu1_M_reg5 (cnu1_f0_M_reg[5]),

        // From the first CNU
        .cnu0_v2c_0 (/*v2c_0*/v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_1 (/*v2c_1*/v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_2 (/*v2c_2*/v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_3 (/*v2c_3*/v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_4 (/*v2c_4*/v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_v2c_5 (/*v2c_5*/v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)]),
        // From the second CNU
        .cnu1_v2c_0 (/*v2c_0*/v2c_latch_0[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_1 (/*v2c_1*/v2c_latch_1[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_2 (/*v2c_2*/v2c_latch_2[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_3 (/*v2c_3*/v2c_latch_3[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_4 (/*v2c_4*/v2c_latch_4[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_v2c_5 (/*v2c_5*/v2c_latch_5[(CNU6_INSTANTIATE_UNIT*j)+1]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset), // offset determing the switch between multi-frame under the following sub-datapath
	
		// Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_0[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_0 (ram_write_dataB_0[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[0])
    );
    // Instantiation of F_1
    wire [QUAN_SIZE-1:0] f1_out[0:3];
    wire [QUAN_SIZE-1:0] cnu0_f1_M_reg [0:CN_DEGREE-1];
    wire [QUAN_SIZE-1:0] cnu1_f1_M_reg [0:CN_DEGREE-1];
    cnu6_f1 u_f1(
		.read_addr_offset_out (read_addr_offset_internal[j][1]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .t_portA (f1_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portB (f1_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        // For the second CNU
        .t_portC (f1_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .t_portD (f1_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the first CNU
        .cnu0_M_reg0 (cnu0_f1_M_reg[0]),
        .cnu0_M_reg1 (cnu0_f1_M_reg[1]),
        .cnu0_M_reg2 (cnu0_f1_M_reg[2]),
        .cnu0_M_reg3 (cnu0_f1_M_reg[3]),
        .cnu0_M_reg4 (cnu0_f1_M_reg[4]),
        .cnu0_M_reg5 (cnu0_f1_M_reg[5]),
        // For the second CNU
        .cnu1_M_reg0 (cnu1_f1_M_reg[0]),
        .cnu1_M_reg1 (cnu1_f1_M_reg[1]),
        .cnu1_M_reg2 (cnu1_f1_M_reg[2]),
        .cnu1_M_reg3 (cnu1_f1_M_reg[3]),
        .cnu1_M_reg4 (cnu1_f1_M_reg[4]),
        .cnu1_M_reg5 (cnu1_f1_M_reg[5]),

        // From the first CNU
        .t_00 (f0_out[0]),
        .t_01 (f0_out[1]),
        .cnu0_v2c_0 (cnu0_f0_M_reg[0]),
        .cnu0_v2c_1 (cnu0_f0_M_reg[1]),
        .cnu0_v2c_2 (cnu0_f0_M_reg[2]),
        .cnu0_v2c_3 (cnu0_f0_M_reg[3]),
        .cnu0_v2c_4 (cnu0_f0_M_reg[4]),
        .cnu0_v2c_5 (cnu0_f0_M_reg[5]),
        // From the second CNU
        .t_02 (f0_out[2]),
        .t_03 (f0_out[3]),
        .cnu1_v2c_0 (cnu1_f0_M_reg[0]),
        .cnu1_v2c_1 (cnu1_f0_M_reg[1]),
        .cnu1_v2c_2 (cnu1_f0_M_reg[2]),
        .cnu1_v2c_3 (cnu1_f0_M_reg[3]),
        .cnu1_v2c_4 (cnu1_f0_M_reg[4]),
        .cnu1_v2c_5 (cnu1_f0_M_reg[5]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset_internal[j][0]), // offset determing the switch between multi-frame under the following sub-datapath

        // Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_1[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_1 (ram_write_dataB_1[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[1])
    );
    // Instantiation of F_2
    wire [QUAN_SIZE-1:0] cnu0_f2_out[0:3];
    wire [QUAN_SIZE-1:0] cnu1_f2_out[0:3];
    wire [QUAN_SIZE-1:0] cnu0_f2_M_reg [0:3];
    wire [QUAN_SIZE-1:0] cnu1_f2_M_reg [0:3];
    cnu6_f2 u_f2(
		.read_addr_offset_out (read_addr_offset_internal[j][2]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .cnu0_t_portA (cnu0_f2_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu0_t_portB (cnu0_f2_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu0_t_portC (cnu0_f2_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu0_t_portD (cnu0_f2_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the second CNU
        .cnu1_t_portA (cnu1_f2_out[0]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu1_t_portB (cnu1_f2_out[1]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu1_t_portC (cnu1_f2_out[2]), // internal signals accounting for each 256-entry partial LUT's output
        .cnu1_t_portD (cnu1_f2_out[3]), // internal signals accounting for each 256-entry partial LUT's output
        // For the first CNU
        .cnu0_M_reg1 (cnu0_f2_M_reg[0]),
        .cnu0_M_reg2 (cnu0_f2_M_reg[1]),
        .cnu0_M_reg4 (cnu0_f2_M_reg[2]),
        .cnu0_M_reg5 (cnu0_f2_M_reg[3]),
        // For the second CNU
        .cnu1_M_reg1 (cnu1_f2_M_reg[0]),
        .cnu1_M_reg2 (cnu1_f2_M_reg[1]),
        .cnu1_M_reg4 (cnu1_f2_M_reg[2]),
        .cnu1_M_reg5 (cnu1_f2_M_reg[3]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset_internal[j][1]), // offset determing the switch between multi-frame under the following sub-datapath

        // From the first CNU
        .t_10 (f1_out[0]),
        .t_11 (f1_out[1]),
        .cnu0_v2c_0 (cnu0_f1_M_reg[0]),
        .cnu0_v2c_1 (cnu0_f1_M_reg[1]),
        .cnu0_v2c_2 (cnu0_f1_M_reg[2]),
        .cnu0_v2c_3 (cnu0_f1_M_reg[3]),
        .cnu0_v2c_4 (cnu0_f1_M_reg[4]),
        .cnu0_v2c_5 (cnu0_f1_M_reg[5]),
        // From the second CNU
        .t_12 (f1_out[2]),
        .t_13 (f1_out[3]),
        .cnu1_v2c_0 (cnu1_f1_M_reg[0]),
        .cnu1_v2c_1 (cnu1_f1_M_reg[1]),
        .cnu1_v2c_2 (cnu1_f1_M_reg[2]),
        .cnu1_v2c_3 (cnu1_f1_M_reg[3]),
        .cnu1_v2c_4 (cnu1_f1_M_reg[4]),
        .cnu1_v2c_5 (cnu1_f1_M_reg[5]),

        // Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_2[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_2 (ram_write_dataB_2[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[2])
    );
    // Instantiation of F_3
    wire [QUAN_SIZE-1:0] cnu0_c2v [0:CN_DEGREE-1];
    wire [QUAN_SIZE-1:0] cnu1_c2v [0:CN_DEGREE-1];
    cnu6_f3 u_f3(
		.read_addr_offset_out (read_addr_offset_outSet[j]), // to forward the current multi-frame offset signal to the next sub-datapath
        // For the first CNU
        .cnu0_c2v_0 (c2v_0[(CNU6_INSTANTIATE_UNIT*j)]), 
        .cnu0_c2v_1 (c2v_1[(CNU6_INSTANTIATE_UNIT*j)]), 
        .cnu0_c2v_2 (c2v_2[(CNU6_INSTANTIATE_UNIT*j)]), 
        .cnu0_c2v_3 (c2v_3[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_c2v_4 (c2v_4[(CNU6_INSTANTIATE_UNIT*j)]),
        .cnu0_c2v_5 (c2v_5[(CNU6_INSTANTIATE_UNIT*j)]), 
        // For the second CNU
        .cnu1_c2v_0 (c2v_0[(CNU6_INSTANTIATE_UNIT*j)+1]), 
        .cnu1_c2v_1 (c2v_1[(CNU6_INSTANTIATE_UNIT*j)+1]), 
        .cnu1_c2v_2 (c2v_2[(CNU6_INSTANTIATE_UNIT*j)+1]), 
        .cnu1_c2v_3 (c2v_3[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_c2v_4 (c2v_4[(CNU6_INSTANTIATE_UNIT*j)+1]),
        .cnu1_c2v_5 (c2v_5[(CNU6_INSTANTIATE_UNIT*j)+1]),

        // From the first CNU
        .cnu0_t_20 (cnu0_f2_out[0]),
        .cnu0_t_21 (cnu0_f2_out[1]),
        .cnu0_t_22 (cnu0_f2_out[2]),
        .cnu0_t_23 (cnu0_f2_out[3]),
        .cnu0_v2c_1 (cnu0_f2_M_reg[0]),
        .cnu0_v2c_2 (cnu0_f2_M_reg[1]),
        .cnu0_v2c_4 (cnu0_f2_M_reg[2]),
        .cnu0_v2c_5 (cnu0_f2_M_reg[3]),
        // From the second CNU
        .cnu1_t_20 (cnu1_f2_out[0]),
        .cnu1_t_21 (cnu1_f2_out[1]),
        .cnu1_t_22 (cnu1_f2_out[2]),
        .cnu1_t_23 (cnu1_f2_out[3]),
        .cnu1_v2c_1 (cnu1_f2_M_reg[0]),
        .cnu1_v2c_2 (cnu1_f2_M_reg[1]),
        .cnu1_v2c_4 (cnu1_f2_M_reg[2]),
        .cnu1_v2c_5 (cnu1_f2_M_reg[3]),

		.read_clk (read_clk),
        .read_addr_offset (read_addr_offset_internal[j][2]), // offset determing the switch between multi-frame under the following sub-datapath

        // Iteration-Update Page Address 
        .page_addr_ram (page_addr_ram_3[CN_PAGE_ADDR_BW+1-1:0]),
        // Iteration-Update Data
        .ram_write_data_3 (ram_write_dataB_3[CN_ROM_RD_BW-1:0]),

        .write_clk (write_clk),
        .ib_ram_we (ib_ram_we[3])
    );
  end
endgenerate

assign c2v_0_out0[QUAN_SIZE-1:0] = c2v_0[0];
assign v2c_0[0] = v2c_0_in0[QUAN_SIZE-1:0];
assign c2v_0_out1[QUAN_SIZE-1:0] = c2v_1[0];
assign v2c_1[0] = v2c_0_in1[QUAN_SIZE-1:0];
assign c2v_0_out2[QUAN_SIZE-1:0] = c2v_2[0];
assign v2c_2[0] = v2c_0_in2[QUAN_SIZE-1:0];
assign c2v_0_out3[QUAN_SIZE-1:0] = c2v_3[0];
assign v2c_3[0] = v2c_0_in3[QUAN_SIZE-1:0];
assign c2v_0_out4[QUAN_SIZE-1:0] = c2v_4[0];
assign v2c_4[0] = v2c_0_in4[QUAN_SIZE-1:0];
assign c2v_0_out5[QUAN_SIZE-1:0] = c2v_5[0];
assign v2c_5[0] = v2c_0_in5[QUAN_SIZE-1:0];
assign c2v_1_out0[QUAN_SIZE-1:0] = c2v_0[1];
assign v2c_0[1] = v2c_1_in0[QUAN_SIZE-1:0];
assign c2v_1_out1[QUAN_SIZE-1:0] = c2v_1[1];
assign v2c_1[1] = v2c_1_in1[QUAN_SIZE-1:0];
assign c2v_1_out2[QUAN_SIZE-1:0] = c2v_2[1];
assign v2c_2[1] = v2c_1_in2[QUAN_SIZE-1:0];
assign c2v_1_out3[QUAN_SIZE-1:0] = c2v_3[1];
assign v2c_3[1] = v2c_1_in3[QUAN_SIZE-1:0];
assign c2v_1_out4[QUAN_SIZE-1:0] = c2v_4[1];
assign v2c_4[1] = v2c_1_in4[QUAN_SIZE-1:0];
assign c2v_1_out5[QUAN_SIZE-1:0] = c2v_5[1];
assign v2c_5[1] = v2c_1_in5[QUAN_SIZE-1:0];
assign c2v_2_out0[QUAN_SIZE-1:0] = c2v_0[2];
assign v2c_0[2] = v2c_2_in0[QUAN_SIZE-1:0];
assign c2v_2_out1[QUAN_SIZE-1:0] = c2v_1[2];
assign v2c_1[2] = v2c_2_in1[QUAN_SIZE-1:0];
assign c2v_2_out2[QUAN_SIZE-1:0] = c2v_2[2];
assign v2c_2[2] = v2c_2_in2[QUAN_SIZE-1:0];
assign c2v_2_out3[QUAN_SIZE-1:0] = c2v_3[2];
assign v2c_3[2] = v2c_2_in3[QUAN_SIZE-1:0];
assign c2v_2_out4[QUAN_SIZE-1:0] = c2v_4[2];
assign v2c_4[2] = v2c_2_in4[QUAN_SIZE-1:0];
assign c2v_2_out5[QUAN_SIZE-1:0] = c2v_5[2];
assign v2c_5[2] = v2c_2_in5[QUAN_SIZE-1:0];
assign c2v_3_out0[QUAN_SIZE-1:0] = c2v_0[3];
assign v2c_0[3] = v2c_3_in0[QUAN_SIZE-1:0];
assign c2v_3_out1[QUAN_SIZE-1:0] = c2v_1[3];
assign v2c_1[3] = v2c_3_in1[QUAN_SIZE-1:0];
assign c2v_3_out2[QUAN_SIZE-1:0] = c2v_2[3];
assign v2c_2[3] = v2c_3_in2[QUAN_SIZE-1:0];
assign c2v_3_out3[QUAN_SIZE-1:0] = c2v_3[3];
assign v2c_3[3] = v2c_3_in3[QUAN_SIZE-1:0];
assign c2v_3_out4[QUAN_SIZE-1:0] = c2v_4[3];
assign v2c_4[3] = v2c_3_in4[QUAN_SIZE-1:0];
assign c2v_3_out5[QUAN_SIZE-1:0] = c2v_5[3];
assign v2c_5[3] = v2c_3_in5[QUAN_SIZE-1:0];
assign c2v_4_out0[QUAN_SIZE-1:0] = c2v_0[4];
assign v2c_0[4] = v2c_4_in0[QUAN_SIZE-1:0];
assign c2v_4_out1[QUAN_SIZE-1:0] = c2v_1[4];
assign v2c_1[4] = v2c_4_in1[QUAN_SIZE-1:0];
assign c2v_4_out2[QUAN_SIZE-1:0] = c2v_2[4];
assign v2c_2[4] = v2c_4_in2[QUAN_SIZE-1:0];
assign c2v_4_out3[QUAN_SIZE-1:0] = c2v_3[4];
assign v2c_3[4] = v2c_4_in3[QUAN_SIZE-1:0];
assign c2v_4_out4[QUAN_SIZE-1:0] = c2v_4[4];
assign v2c_4[4] = v2c_4_in4[QUAN_SIZE-1:0];
assign c2v_4_out5[QUAN_SIZE-1:0] = c2v_5[4];
assign v2c_5[4] = v2c_4_in5[QUAN_SIZE-1:0];
assign c2v_5_out0[QUAN_SIZE-1:0] = c2v_0[5];
assign v2c_0[5] = v2c_5_in0[QUAN_SIZE-1:0];
assign c2v_5_out1[QUAN_SIZE-1:0] = c2v_1[5];
assign v2c_1[5] = v2c_5_in1[QUAN_SIZE-1:0];
assign c2v_5_out2[QUAN_SIZE-1:0] = c2v_2[5];
assign v2c_2[5] = v2c_5_in2[QUAN_SIZE-1:0];
assign c2v_5_out3[QUAN_SIZE-1:0] = c2v_3[5];
assign v2c_3[5] = v2c_5_in3[QUAN_SIZE-1:0];
assign c2v_5_out4[QUAN_SIZE-1:0] = c2v_4[5];
assign v2c_4[5] = v2c_5_in4[QUAN_SIZE-1:0];
assign c2v_5_out5[QUAN_SIZE-1:0] = c2v_5[5];
assign v2c_5[5] = v2c_5_in5[QUAN_SIZE-1:0];
assign c2v_6_out0[QUAN_SIZE-1:0] = c2v_0[6];
assign v2c_0[6] = v2c_6_in0[QUAN_SIZE-1:0];
assign c2v_6_out1[QUAN_SIZE-1:0] = c2v_1[6];
assign v2c_1[6] = v2c_6_in1[QUAN_SIZE-1:0];
assign c2v_6_out2[QUAN_SIZE-1:0] = c2v_2[6];
assign v2c_2[6] = v2c_6_in2[QUAN_SIZE-1:0];
assign c2v_6_out3[QUAN_SIZE-1:0] = c2v_3[6];
assign v2c_3[6] = v2c_6_in3[QUAN_SIZE-1:0];
assign c2v_6_out4[QUAN_SIZE-1:0] = c2v_4[6];
assign v2c_4[6] = v2c_6_in4[QUAN_SIZE-1:0];
assign c2v_6_out5[QUAN_SIZE-1:0] = c2v_5[6];
assign v2c_5[6] = v2c_6_in5[QUAN_SIZE-1:0];
assign c2v_7_out0[QUAN_SIZE-1:0] = c2v_0[7];
assign v2c_0[7] = v2c_7_in0[QUAN_SIZE-1:0];
assign c2v_7_out1[QUAN_SIZE-1:0] = c2v_1[7];
assign v2c_1[7] = v2c_7_in1[QUAN_SIZE-1:0];
assign c2v_7_out2[QUAN_SIZE-1:0] = c2v_2[7];
assign v2c_2[7] = v2c_7_in2[QUAN_SIZE-1:0];
assign c2v_7_out3[QUAN_SIZE-1:0] = c2v_3[7];
assign v2c_3[7] = v2c_7_in3[QUAN_SIZE-1:0];
assign c2v_7_out4[QUAN_SIZE-1:0] = c2v_4[7];
assign v2c_4[7] = v2c_7_in4[QUAN_SIZE-1:0];
assign c2v_7_out5[QUAN_SIZE-1:0] = c2v_5[7];
assign v2c_5[7] = v2c_7_in5[QUAN_SIZE-1:0];
assign c2v_8_out0[QUAN_SIZE-1:0] = c2v_0[8];
assign v2c_0[8] = v2c_8_in0[QUAN_SIZE-1:0];
assign c2v_8_out1[QUAN_SIZE-1:0] = c2v_1[8];
assign v2c_1[8] = v2c_8_in1[QUAN_SIZE-1:0];
assign c2v_8_out2[QUAN_SIZE-1:0] = c2v_2[8];
assign v2c_2[8] = v2c_8_in2[QUAN_SIZE-1:0];
assign c2v_8_out3[QUAN_SIZE-1:0] = c2v_3[8];
assign v2c_3[8] = v2c_8_in3[QUAN_SIZE-1:0];
assign c2v_8_out4[QUAN_SIZE-1:0] = c2v_4[8];
assign v2c_4[8] = v2c_8_in4[QUAN_SIZE-1:0];
assign c2v_8_out5[QUAN_SIZE-1:0] = c2v_5[8];
assign v2c_5[8] = v2c_8_in5[QUAN_SIZE-1:0];
assign c2v_9_out0[QUAN_SIZE-1:0] = c2v_0[9];
assign v2c_0[9] = v2c_9_in0[QUAN_SIZE-1:0];
assign c2v_9_out1[QUAN_SIZE-1:0] = c2v_1[9];
assign v2c_1[9] = v2c_9_in1[QUAN_SIZE-1:0];
assign c2v_9_out2[QUAN_SIZE-1:0] = c2v_2[9];
assign v2c_2[9] = v2c_9_in2[QUAN_SIZE-1:0];
assign c2v_9_out3[QUAN_SIZE-1:0] = c2v_3[9];
assign v2c_3[9] = v2c_9_in3[QUAN_SIZE-1:0];
assign c2v_9_out4[QUAN_SIZE-1:0] = c2v_4[9];
assign v2c_4[9] = v2c_9_in4[QUAN_SIZE-1:0];
assign c2v_9_out5[QUAN_SIZE-1:0] = c2v_5[9];
assign v2c_5[9] = v2c_9_in5[QUAN_SIZE-1:0];
assign c2v_10_out0[QUAN_SIZE-1:0] = c2v_0[10];
assign v2c_0[10] = v2c_10_in0[QUAN_SIZE-1:0];
assign c2v_10_out1[QUAN_SIZE-1:0] = c2v_1[10];
assign v2c_1[10] = v2c_10_in1[QUAN_SIZE-1:0];
assign c2v_10_out2[QUAN_SIZE-1:0] = c2v_2[10];
assign v2c_2[10] = v2c_10_in2[QUAN_SIZE-1:0];
assign c2v_10_out3[QUAN_SIZE-1:0] = c2v_3[10];
assign v2c_3[10] = v2c_10_in3[QUAN_SIZE-1:0];
assign c2v_10_out4[QUAN_SIZE-1:0] = c2v_4[10];
assign v2c_4[10] = v2c_10_in4[QUAN_SIZE-1:0];
assign c2v_10_out5[QUAN_SIZE-1:0] = c2v_5[10];
assign v2c_5[10] = v2c_10_in5[QUAN_SIZE-1:0];
assign c2v_11_out0[QUAN_SIZE-1:0] = c2v_0[11];
assign v2c_0[11] = v2c_11_in0[QUAN_SIZE-1:0];
assign c2v_11_out1[QUAN_SIZE-1:0] = c2v_1[11];
assign v2c_1[11] = v2c_11_in1[QUAN_SIZE-1:0];
assign c2v_11_out2[QUAN_SIZE-1:0] = c2v_2[11];
assign v2c_2[11] = v2c_11_in2[QUAN_SIZE-1:0];
assign c2v_11_out3[QUAN_SIZE-1:0] = c2v_3[11];
assign v2c_3[11] = v2c_11_in3[QUAN_SIZE-1:0];
assign c2v_11_out4[QUAN_SIZE-1:0] = c2v_4[11];
assign v2c_4[11] = v2c_11_in4[QUAN_SIZE-1:0];
assign c2v_11_out5[QUAN_SIZE-1:0] = c2v_5[11];
assign v2c_5[11] = v2c_11_in5[QUAN_SIZE-1:0];
assign c2v_12_out0[QUAN_SIZE-1:0] = c2v_0[12];
assign v2c_0[12] = v2c_12_in0[QUAN_SIZE-1:0];
assign c2v_12_out1[QUAN_SIZE-1:0] = c2v_1[12];
assign v2c_1[12] = v2c_12_in1[QUAN_SIZE-1:0];
assign c2v_12_out2[QUAN_SIZE-1:0] = c2v_2[12];
assign v2c_2[12] = v2c_12_in2[QUAN_SIZE-1:0];
assign c2v_12_out3[QUAN_SIZE-1:0] = c2v_3[12];
assign v2c_3[12] = v2c_12_in3[QUAN_SIZE-1:0];
assign c2v_12_out4[QUAN_SIZE-1:0] = c2v_4[12];
assign v2c_4[12] = v2c_12_in4[QUAN_SIZE-1:0];
assign c2v_12_out5[QUAN_SIZE-1:0] = c2v_5[12];
assign v2c_5[12] = v2c_12_in5[QUAN_SIZE-1:0];
assign c2v_13_out0[QUAN_SIZE-1:0] = c2v_0[13];
assign v2c_0[13] = v2c_13_in0[QUAN_SIZE-1:0];
assign c2v_13_out1[QUAN_SIZE-1:0] = c2v_1[13];
assign v2c_1[13] = v2c_13_in1[QUAN_SIZE-1:0];
assign c2v_13_out2[QUAN_SIZE-1:0] = c2v_2[13];
assign v2c_2[13] = v2c_13_in2[QUAN_SIZE-1:0];
assign c2v_13_out3[QUAN_SIZE-1:0] = c2v_3[13];
assign v2c_3[13] = v2c_13_in3[QUAN_SIZE-1:0];
assign c2v_13_out4[QUAN_SIZE-1:0] = c2v_4[13];
assign v2c_4[13] = v2c_13_in4[QUAN_SIZE-1:0];
assign c2v_13_out5[QUAN_SIZE-1:0] = c2v_5[13];
assign v2c_5[13] = v2c_13_in5[QUAN_SIZE-1:0];
assign c2v_14_out0[QUAN_SIZE-1:0] = c2v_0[14];
assign v2c_0[14] = v2c_14_in0[QUAN_SIZE-1:0];
assign c2v_14_out1[QUAN_SIZE-1:0] = c2v_1[14];
assign v2c_1[14] = v2c_14_in1[QUAN_SIZE-1:0];
assign c2v_14_out2[QUAN_SIZE-1:0] = c2v_2[14];
assign v2c_2[14] = v2c_14_in2[QUAN_SIZE-1:0];
assign c2v_14_out3[QUAN_SIZE-1:0] = c2v_3[14];
assign v2c_3[14] = v2c_14_in3[QUAN_SIZE-1:0];
assign c2v_14_out4[QUAN_SIZE-1:0] = c2v_4[14];
assign v2c_4[14] = v2c_14_in4[QUAN_SIZE-1:0];
assign c2v_14_out5[QUAN_SIZE-1:0] = c2v_5[14];
assign v2c_5[14] = v2c_14_in5[QUAN_SIZE-1:0];
assign c2v_15_out0[QUAN_SIZE-1:0] = c2v_0[15];
assign v2c_0[15] = v2c_15_in0[QUAN_SIZE-1:0];
assign c2v_15_out1[QUAN_SIZE-1:0] = c2v_1[15];
assign v2c_1[15] = v2c_15_in1[QUAN_SIZE-1:0];
assign c2v_15_out2[QUAN_SIZE-1:0] = c2v_2[15];
assign v2c_2[15] = v2c_15_in2[QUAN_SIZE-1:0];
assign c2v_15_out3[QUAN_SIZE-1:0] = c2v_3[15];
assign v2c_3[15] = v2c_15_in3[QUAN_SIZE-1:0];
assign c2v_15_out4[QUAN_SIZE-1:0] = c2v_4[15];
assign v2c_4[15] = v2c_15_in4[QUAN_SIZE-1:0];
assign c2v_15_out5[QUAN_SIZE-1:0] = c2v_5[15];
assign v2c_5[15] = v2c_15_in5[QUAN_SIZE-1:0];
assign c2v_16_out0[QUAN_SIZE-1:0] = c2v_0[16];
assign v2c_0[16] = v2c_16_in0[QUAN_SIZE-1:0];
assign c2v_16_out1[QUAN_SIZE-1:0] = c2v_1[16];
assign v2c_1[16] = v2c_16_in1[QUAN_SIZE-1:0];
assign c2v_16_out2[QUAN_SIZE-1:0] = c2v_2[16];
assign v2c_2[16] = v2c_16_in2[QUAN_SIZE-1:0];
assign c2v_16_out3[QUAN_SIZE-1:0] = c2v_3[16];
assign v2c_3[16] = v2c_16_in3[QUAN_SIZE-1:0];
assign c2v_16_out4[QUAN_SIZE-1:0] = c2v_4[16];
assign v2c_4[16] = v2c_16_in4[QUAN_SIZE-1:0];
assign c2v_16_out5[QUAN_SIZE-1:0] = c2v_5[16];
assign v2c_5[16] = v2c_16_in5[QUAN_SIZE-1:0];
assign c2v_17_out0[QUAN_SIZE-1:0] = c2v_0[17];
assign v2c_0[17] = v2c_17_in0[QUAN_SIZE-1:0];
assign c2v_17_out1[QUAN_SIZE-1:0] = c2v_1[17];
assign v2c_1[17] = v2c_17_in1[QUAN_SIZE-1:0];
assign c2v_17_out2[QUAN_SIZE-1:0] = c2v_2[17];
assign v2c_2[17] = v2c_17_in2[QUAN_SIZE-1:0];
assign c2v_17_out3[QUAN_SIZE-1:0] = c2v_3[17];
assign v2c_3[17] = v2c_17_in3[QUAN_SIZE-1:0];
assign c2v_17_out4[QUAN_SIZE-1:0] = c2v_4[17];
assign v2c_4[17] = v2c_17_in4[QUAN_SIZE-1:0];
assign c2v_17_out5[QUAN_SIZE-1:0] = c2v_5[17];
assign v2c_5[17] = v2c_17_in5[QUAN_SIZE-1:0];
assign c2v_18_out0[QUAN_SIZE-1:0] = c2v_0[18];
assign v2c_0[18] = v2c_18_in0[QUAN_SIZE-1:0];
assign c2v_18_out1[QUAN_SIZE-1:0] = c2v_1[18];
assign v2c_1[18] = v2c_18_in1[QUAN_SIZE-1:0];
assign c2v_18_out2[QUAN_SIZE-1:0] = c2v_2[18];
assign v2c_2[18] = v2c_18_in2[QUAN_SIZE-1:0];
assign c2v_18_out3[QUAN_SIZE-1:0] = c2v_3[18];
assign v2c_3[18] = v2c_18_in3[QUAN_SIZE-1:0];
assign c2v_18_out4[QUAN_SIZE-1:0] = c2v_4[18];
assign v2c_4[18] = v2c_18_in4[QUAN_SIZE-1:0];
assign c2v_18_out5[QUAN_SIZE-1:0] = c2v_5[18];
assign v2c_5[18] = v2c_18_in5[QUAN_SIZE-1:0];
assign c2v_19_out0[QUAN_SIZE-1:0] = c2v_0[19];
assign v2c_0[19] = v2c_19_in0[QUAN_SIZE-1:0];
assign c2v_19_out1[QUAN_SIZE-1:0] = c2v_1[19];
assign v2c_1[19] = v2c_19_in1[QUAN_SIZE-1:0];
assign c2v_19_out2[QUAN_SIZE-1:0] = c2v_2[19];
assign v2c_2[19] = v2c_19_in2[QUAN_SIZE-1:0];
assign c2v_19_out3[QUAN_SIZE-1:0] = c2v_3[19];
assign v2c_3[19] = v2c_19_in3[QUAN_SIZE-1:0];
assign c2v_19_out4[QUAN_SIZE-1:0] = c2v_4[19];
assign v2c_4[19] = v2c_19_in4[QUAN_SIZE-1:0];
assign c2v_19_out5[QUAN_SIZE-1:0] = c2v_5[19];
assign v2c_5[19] = v2c_19_in5[QUAN_SIZE-1:0];
assign c2v_20_out0[QUAN_SIZE-1:0] = c2v_0[20];
assign v2c_0[20] = v2c_20_in0[QUAN_SIZE-1:0];
assign c2v_20_out1[QUAN_SIZE-1:0] = c2v_1[20];
assign v2c_1[20] = v2c_20_in1[QUAN_SIZE-1:0];
assign c2v_20_out2[QUAN_SIZE-1:0] = c2v_2[20];
assign v2c_2[20] = v2c_20_in2[QUAN_SIZE-1:0];
assign c2v_20_out3[QUAN_SIZE-1:0] = c2v_3[20];
assign v2c_3[20] = v2c_20_in3[QUAN_SIZE-1:0];
assign c2v_20_out4[QUAN_SIZE-1:0] = c2v_4[20];
assign v2c_4[20] = v2c_20_in4[QUAN_SIZE-1:0];
assign c2v_20_out5[QUAN_SIZE-1:0] = c2v_5[20];
assign v2c_5[20] = v2c_20_in5[QUAN_SIZE-1:0];
assign c2v_21_out0[QUAN_SIZE-1:0] = c2v_0[21];
assign v2c_0[21] = v2c_21_in0[QUAN_SIZE-1:0];
assign c2v_21_out1[QUAN_SIZE-1:0] = c2v_1[21];
assign v2c_1[21] = v2c_21_in1[QUAN_SIZE-1:0];
assign c2v_21_out2[QUAN_SIZE-1:0] = c2v_2[21];
assign v2c_2[21] = v2c_21_in2[QUAN_SIZE-1:0];
assign c2v_21_out3[QUAN_SIZE-1:0] = c2v_3[21];
assign v2c_3[21] = v2c_21_in3[QUAN_SIZE-1:0];
assign c2v_21_out4[QUAN_SIZE-1:0] = c2v_4[21];
assign v2c_4[21] = v2c_21_in4[QUAN_SIZE-1:0];
assign c2v_21_out5[QUAN_SIZE-1:0] = c2v_5[21];
assign v2c_5[21] = v2c_21_in5[QUAN_SIZE-1:0];
assign c2v_22_out0[QUAN_SIZE-1:0] = c2v_0[22];
assign v2c_0[22] = v2c_22_in0[QUAN_SIZE-1:0];
assign c2v_22_out1[QUAN_SIZE-1:0] = c2v_1[22];
assign v2c_1[22] = v2c_22_in1[QUAN_SIZE-1:0];
assign c2v_22_out2[QUAN_SIZE-1:0] = c2v_2[22];
assign v2c_2[22] = v2c_22_in2[QUAN_SIZE-1:0];
assign c2v_22_out3[QUAN_SIZE-1:0] = c2v_3[22];
assign v2c_3[22] = v2c_22_in3[QUAN_SIZE-1:0];
assign c2v_22_out4[QUAN_SIZE-1:0] = c2v_4[22];
assign v2c_4[22] = v2c_22_in4[QUAN_SIZE-1:0];
assign c2v_22_out5[QUAN_SIZE-1:0] = c2v_5[22];
assign v2c_5[22] = v2c_22_in5[QUAN_SIZE-1:0];
assign c2v_23_out0[QUAN_SIZE-1:0] = c2v_0[23];
assign v2c_0[23] = v2c_23_in0[QUAN_SIZE-1:0];
assign c2v_23_out1[QUAN_SIZE-1:0] = c2v_1[23];
assign v2c_1[23] = v2c_23_in1[QUAN_SIZE-1:0];
assign c2v_23_out2[QUAN_SIZE-1:0] = c2v_2[23];
assign v2c_2[23] = v2c_23_in2[QUAN_SIZE-1:0];
assign c2v_23_out3[QUAN_SIZE-1:0] = c2v_3[23];
assign v2c_3[23] = v2c_23_in3[QUAN_SIZE-1:0];
assign c2v_23_out4[QUAN_SIZE-1:0] = c2v_4[23];
assign v2c_4[23] = v2c_23_in4[QUAN_SIZE-1:0];
assign c2v_23_out5[QUAN_SIZE-1:0] = c2v_5[23];
assign v2c_5[23] = v2c_23_in5[QUAN_SIZE-1:0];
assign c2v_24_out0[QUAN_SIZE-1:0] = c2v_0[24];
assign v2c_0[24] = v2c_24_in0[QUAN_SIZE-1:0];
assign c2v_24_out1[QUAN_SIZE-1:0] = c2v_1[24];
assign v2c_1[24] = v2c_24_in1[QUAN_SIZE-1:0];
assign c2v_24_out2[QUAN_SIZE-1:0] = c2v_2[24];
assign v2c_2[24] = v2c_24_in2[QUAN_SIZE-1:0];
assign c2v_24_out3[QUAN_SIZE-1:0] = c2v_3[24];
assign v2c_3[24] = v2c_24_in3[QUAN_SIZE-1:0];
assign c2v_24_out4[QUAN_SIZE-1:0] = c2v_4[24];
assign v2c_4[24] = v2c_24_in4[QUAN_SIZE-1:0];
assign c2v_24_out5[QUAN_SIZE-1:0] = c2v_5[24];
assign v2c_5[24] = v2c_24_in5[QUAN_SIZE-1:0];
assign c2v_25_out0[QUAN_SIZE-1:0] = c2v_0[25];
assign v2c_0[25] = v2c_25_in0[QUAN_SIZE-1:0];
assign c2v_25_out1[QUAN_SIZE-1:0] = c2v_1[25];
assign v2c_1[25] = v2c_25_in1[QUAN_SIZE-1:0];
assign c2v_25_out2[QUAN_SIZE-1:0] = c2v_2[25];
assign v2c_2[25] = v2c_25_in2[QUAN_SIZE-1:0];
assign c2v_25_out3[QUAN_SIZE-1:0] = c2v_3[25];
assign v2c_3[25] = v2c_25_in3[QUAN_SIZE-1:0];
assign c2v_25_out4[QUAN_SIZE-1:0] = c2v_4[25];
assign v2c_4[25] = v2c_25_in4[QUAN_SIZE-1:0];
assign c2v_25_out5[QUAN_SIZE-1:0] = c2v_5[25];
assign v2c_5[25] = v2c_25_in5[QUAN_SIZE-1:0];
assign c2v_26_out0[QUAN_SIZE-1:0] = c2v_0[26];
assign v2c_0[26] = v2c_26_in0[QUAN_SIZE-1:0];
assign c2v_26_out1[QUAN_SIZE-1:0] = c2v_1[26];
assign v2c_1[26] = v2c_26_in1[QUAN_SIZE-1:0];
assign c2v_26_out2[QUAN_SIZE-1:0] = c2v_2[26];
assign v2c_2[26] = v2c_26_in2[QUAN_SIZE-1:0];
assign c2v_26_out3[QUAN_SIZE-1:0] = c2v_3[26];
assign v2c_3[26] = v2c_26_in3[QUAN_SIZE-1:0];
assign c2v_26_out4[QUAN_SIZE-1:0] = c2v_4[26];
assign v2c_4[26] = v2c_26_in4[QUAN_SIZE-1:0];
assign c2v_26_out5[QUAN_SIZE-1:0] = c2v_5[26];
assign v2c_5[26] = v2c_26_in5[QUAN_SIZE-1:0];
assign c2v_27_out0[QUAN_SIZE-1:0] = c2v_0[27];
assign v2c_0[27] = v2c_27_in0[QUAN_SIZE-1:0];
assign c2v_27_out1[QUAN_SIZE-1:0] = c2v_1[27];
assign v2c_1[27] = v2c_27_in1[QUAN_SIZE-1:0];
assign c2v_27_out2[QUAN_SIZE-1:0] = c2v_2[27];
assign v2c_2[27] = v2c_27_in2[QUAN_SIZE-1:0];
assign c2v_27_out3[QUAN_SIZE-1:0] = c2v_3[27];
assign v2c_3[27] = v2c_27_in3[QUAN_SIZE-1:0];
assign c2v_27_out4[QUAN_SIZE-1:0] = c2v_4[27];
assign v2c_4[27] = v2c_27_in4[QUAN_SIZE-1:0];
assign c2v_27_out5[QUAN_SIZE-1:0] = c2v_5[27];
assign v2c_5[27] = v2c_27_in5[QUAN_SIZE-1:0];
assign c2v_28_out0[QUAN_SIZE-1:0] = c2v_0[28];
assign v2c_0[28] = v2c_28_in0[QUAN_SIZE-1:0];
assign c2v_28_out1[QUAN_SIZE-1:0] = c2v_1[28];
assign v2c_1[28] = v2c_28_in1[QUAN_SIZE-1:0];
assign c2v_28_out2[QUAN_SIZE-1:0] = c2v_2[28];
assign v2c_2[28] = v2c_28_in2[QUAN_SIZE-1:0];
assign c2v_28_out3[QUAN_SIZE-1:0] = c2v_3[28];
assign v2c_3[28] = v2c_28_in3[QUAN_SIZE-1:0];
assign c2v_28_out4[QUAN_SIZE-1:0] = c2v_4[28];
assign v2c_4[28] = v2c_28_in4[QUAN_SIZE-1:0];
assign c2v_28_out5[QUAN_SIZE-1:0] = c2v_5[28];
assign v2c_5[28] = v2c_28_in5[QUAN_SIZE-1:0];
assign c2v_29_out0[QUAN_SIZE-1:0] = c2v_0[29];
assign v2c_0[29] = v2c_29_in0[QUAN_SIZE-1:0];
assign c2v_29_out1[QUAN_SIZE-1:0] = c2v_1[29];
assign v2c_1[29] = v2c_29_in1[QUAN_SIZE-1:0];
assign c2v_29_out2[QUAN_SIZE-1:0] = c2v_2[29];
assign v2c_2[29] = v2c_29_in2[QUAN_SIZE-1:0];
assign c2v_29_out3[QUAN_SIZE-1:0] = c2v_3[29];
assign v2c_3[29] = v2c_29_in3[QUAN_SIZE-1:0];
assign c2v_29_out4[QUAN_SIZE-1:0] = c2v_4[29];
assign v2c_4[29] = v2c_29_in4[QUAN_SIZE-1:0];
assign c2v_29_out5[QUAN_SIZE-1:0] = c2v_5[29];
assign v2c_5[29] = v2c_29_in5[QUAN_SIZE-1:0];
assign c2v_30_out0[QUAN_SIZE-1:0] = c2v_0[30];
assign v2c_0[30] = v2c_30_in0[QUAN_SIZE-1:0];
assign c2v_30_out1[QUAN_SIZE-1:0] = c2v_1[30];
assign v2c_1[30] = v2c_30_in1[QUAN_SIZE-1:0];
assign c2v_30_out2[QUAN_SIZE-1:0] = c2v_2[30];
assign v2c_2[30] = v2c_30_in2[QUAN_SIZE-1:0];
assign c2v_30_out3[QUAN_SIZE-1:0] = c2v_3[30];
assign v2c_3[30] = v2c_30_in3[QUAN_SIZE-1:0];
assign c2v_30_out4[QUAN_SIZE-1:0] = c2v_4[30];
assign v2c_4[30] = v2c_30_in4[QUAN_SIZE-1:0];
assign c2v_30_out5[QUAN_SIZE-1:0] = c2v_5[30];
assign v2c_5[30] = v2c_30_in5[QUAN_SIZE-1:0];
assign c2v_31_out0[QUAN_SIZE-1:0] = c2v_0[31];
assign v2c_0[31] = v2c_31_in0[QUAN_SIZE-1:0];
assign c2v_31_out1[QUAN_SIZE-1:0] = c2v_1[31];
assign v2c_1[31] = v2c_31_in1[QUAN_SIZE-1:0];
assign c2v_31_out2[QUAN_SIZE-1:0] = c2v_2[31];
assign v2c_2[31] = v2c_31_in2[QUAN_SIZE-1:0];
assign c2v_31_out3[QUAN_SIZE-1:0] = c2v_3[31];
assign v2c_3[31] = v2c_31_in3[QUAN_SIZE-1:0];
assign c2v_31_out4[QUAN_SIZE-1:0] = c2v_4[31];
assign v2c_4[31] = v2c_31_in4[QUAN_SIZE-1:0];
assign c2v_31_out5[QUAN_SIZE-1:0] = c2v_5[31];
assign v2c_5[31] = v2c_31_in5[QUAN_SIZE-1:0];
assign c2v_32_out0[QUAN_SIZE-1:0] = c2v_0[32];
assign v2c_0[32] = v2c_32_in0[QUAN_SIZE-1:0];
assign c2v_32_out1[QUAN_SIZE-1:0] = c2v_1[32];
assign v2c_1[32] = v2c_32_in1[QUAN_SIZE-1:0];
assign c2v_32_out2[QUAN_SIZE-1:0] = c2v_2[32];
assign v2c_2[32] = v2c_32_in2[QUAN_SIZE-1:0];
assign c2v_32_out3[QUAN_SIZE-1:0] = c2v_3[32];
assign v2c_3[32] = v2c_32_in3[QUAN_SIZE-1:0];
assign c2v_32_out4[QUAN_SIZE-1:0] = c2v_4[32];
assign v2c_4[32] = v2c_32_in4[QUAN_SIZE-1:0];
assign c2v_32_out5[QUAN_SIZE-1:0] = c2v_5[32];
assign v2c_5[32] = v2c_32_in5[QUAN_SIZE-1:0];
assign c2v_33_out0[QUAN_SIZE-1:0] = c2v_0[33];
assign v2c_0[33] = v2c_33_in0[QUAN_SIZE-1:0];
assign c2v_33_out1[QUAN_SIZE-1:0] = c2v_1[33];
assign v2c_1[33] = v2c_33_in1[QUAN_SIZE-1:0];
assign c2v_33_out2[QUAN_SIZE-1:0] = c2v_2[33];
assign v2c_2[33] = v2c_33_in2[QUAN_SIZE-1:0];
assign c2v_33_out3[QUAN_SIZE-1:0] = c2v_3[33];
assign v2c_3[33] = v2c_33_in3[QUAN_SIZE-1:0];
assign c2v_33_out4[QUAN_SIZE-1:0] = c2v_4[33];
assign v2c_4[33] = v2c_33_in4[QUAN_SIZE-1:0];
assign c2v_33_out5[QUAN_SIZE-1:0] = c2v_5[33];
assign v2c_5[33] = v2c_33_in5[QUAN_SIZE-1:0];
assign c2v_34_out0[QUAN_SIZE-1:0] = c2v_0[34];
assign v2c_0[34] = v2c_34_in0[QUAN_SIZE-1:0];
assign c2v_34_out1[QUAN_SIZE-1:0] = c2v_1[34];
assign v2c_1[34] = v2c_34_in1[QUAN_SIZE-1:0];
assign c2v_34_out2[QUAN_SIZE-1:0] = c2v_2[34];
assign v2c_2[34] = v2c_34_in2[QUAN_SIZE-1:0];
assign c2v_34_out3[QUAN_SIZE-1:0] = c2v_3[34];
assign v2c_3[34] = v2c_34_in3[QUAN_SIZE-1:0];
assign c2v_34_out4[QUAN_SIZE-1:0] = c2v_4[34];
assign v2c_4[34] = v2c_34_in4[QUAN_SIZE-1:0];
assign c2v_34_out5[QUAN_SIZE-1:0] = c2v_5[34];
assign v2c_5[34] = v2c_34_in5[QUAN_SIZE-1:0];
assign c2v_35_out0[QUAN_SIZE-1:0] = c2v_0[35];
assign v2c_0[35] = v2c_35_in0[QUAN_SIZE-1:0];
assign c2v_35_out1[QUAN_SIZE-1:0] = c2v_1[35];
assign v2c_1[35] = v2c_35_in1[QUAN_SIZE-1:0];
assign c2v_35_out2[QUAN_SIZE-1:0] = c2v_2[35];
assign v2c_2[35] = v2c_35_in2[QUAN_SIZE-1:0];
assign c2v_35_out3[QUAN_SIZE-1:0] = c2v_3[35];
assign v2c_3[35] = v2c_35_in3[QUAN_SIZE-1:0];
assign c2v_35_out4[QUAN_SIZE-1:0] = c2v_4[35];
assign v2c_4[35] = v2c_35_in4[QUAN_SIZE-1:0];
assign c2v_35_out5[QUAN_SIZE-1:0] = c2v_5[35];
assign v2c_5[35] = v2c_35_in5[QUAN_SIZE-1:0];
assign c2v_36_out0[QUAN_SIZE-1:0] = c2v_0[36];
assign v2c_0[36] = v2c_36_in0[QUAN_SIZE-1:0];
assign c2v_36_out1[QUAN_SIZE-1:0] = c2v_1[36];
assign v2c_1[36] = v2c_36_in1[QUAN_SIZE-1:0];
assign c2v_36_out2[QUAN_SIZE-1:0] = c2v_2[36];
assign v2c_2[36] = v2c_36_in2[QUAN_SIZE-1:0];
assign c2v_36_out3[QUAN_SIZE-1:0] = c2v_3[36];
assign v2c_3[36] = v2c_36_in3[QUAN_SIZE-1:0];
assign c2v_36_out4[QUAN_SIZE-1:0] = c2v_4[36];
assign v2c_4[36] = v2c_36_in4[QUAN_SIZE-1:0];
assign c2v_36_out5[QUAN_SIZE-1:0] = c2v_5[36];
assign v2c_5[36] = v2c_36_in5[QUAN_SIZE-1:0];
assign c2v_37_out0[QUAN_SIZE-1:0] = c2v_0[37];
assign v2c_0[37] = v2c_37_in0[QUAN_SIZE-1:0];
assign c2v_37_out1[QUAN_SIZE-1:0] = c2v_1[37];
assign v2c_1[37] = v2c_37_in1[QUAN_SIZE-1:0];
assign c2v_37_out2[QUAN_SIZE-1:0] = c2v_2[37];
assign v2c_2[37] = v2c_37_in2[QUAN_SIZE-1:0];
assign c2v_37_out3[QUAN_SIZE-1:0] = c2v_3[37];
assign v2c_3[37] = v2c_37_in3[QUAN_SIZE-1:0];
assign c2v_37_out4[QUAN_SIZE-1:0] = c2v_4[37];
assign v2c_4[37] = v2c_37_in4[QUAN_SIZE-1:0];
assign c2v_37_out5[QUAN_SIZE-1:0] = c2v_5[37];
assign v2c_5[37] = v2c_37_in5[QUAN_SIZE-1:0];
assign c2v_38_out0[QUAN_SIZE-1:0] = c2v_0[38];
assign v2c_0[38] = v2c_38_in0[QUAN_SIZE-1:0];
assign c2v_38_out1[QUAN_SIZE-1:0] = c2v_1[38];
assign v2c_1[38] = v2c_38_in1[QUAN_SIZE-1:0];
assign c2v_38_out2[QUAN_SIZE-1:0] = c2v_2[38];
assign v2c_2[38] = v2c_38_in2[QUAN_SIZE-1:0];
assign c2v_38_out3[QUAN_SIZE-1:0] = c2v_3[38];
assign v2c_3[38] = v2c_38_in3[QUAN_SIZE-1:0];
assign c2v_38_out4[QUAN_SIZE-1:0] = c2v_4[38];
assign v2c_4[38] = v2c_38_in4[QUAN_SIZE-1:0];
assign c2v_38_out5[QUAN_SIZE-1:0] = c2v_5[38];
assign v2c_5[38] = v2c_38_in5[QUAN_SIZE-1:0];
assign c2v_39_out0[QUAN_SIZE-1:0] = c2v_0[39];
assign v2c_0[39] = v2c_39_in0[QUAN_SIZE-1:0];
assign c2v_39_out1[QUAN_SIZE-1:0] = c2v_1[39];
assign v2c_1[39] = v2c_39_in1[QUAN_SIZE-1:0];
assign c2v_39_out2[QUAN_SIZE-1:0] = c2v_2[39];
assign v2c_2[39] = v2c_39_in2[QUAN_SIZE-1:0];
assign c2v_39_out3[QUAN_SIZE-1:0] = c2v_3[39];
assign v2c_3[39] = v2c_39_in3[QUAN_SIZE-1:0];
assign c2v_39_out4[QUAN_SIZE-1:0] = c2v_4[39];
assign v2c_4[39] = v2c_39_in4[QUAN_SIZE-1:0];
assign c2v_39_out5[QUAN_SIZE-1:0] = c2v_5[39];
assign v2c_5[39] = v2c_39_in5[QUAN_SIZE-1:0];
assign c2v_40_out0[QUAN_SIZE-1:0] = c2v_0[40];
assign v2c_0[40] = v2c_40_in0[QUAN_SIZE-1:0];
assign c2v_40_out1[QUAN_SIZE-1:0] = c2v_1[40];
assign v2c_1[40] = v2c_40_in1[QUAN_SIZE-1:0];
assign c2v_40_out2[QUAN_SIZE-1:0] = c2v_2[40];
assign v2c_2[40] = v2c_40_in2[QUAN_SIZE-1:0];
assign c2v_40_out3[QUAN_SIZE-1:0] = c2v_3[40];
assign v2c_3[40] = v2c_40_in3[QUAN_SIZE-1:0];
assign c2v_40_out4[QUAN_SIZE-1:0] = c2v_4[40];
assign v2c_4[40] = v2c_40_in4[QUAN_SIZE-1:0];
assign c2v_40_out5[QUAN_SIZE-1:0] = c2v_5[40];
assign v2c_5[40] = v2c_40_in5[QUAN_SIZE-1:0];
assign c2v_41_out0[QUAN_SIZE-1:0] = c2v_0[41];
assign v2c_0[41] = v2c_41_in0[QUAN_SIZE-1:0];
assign c2v_41_out1[QUAN_SIZE-1:0] = c2v_1[41];
assign v2c_1[41] = v2c_41_in1[QUAN_SIZE-1:0];
assign c2v_41_out2[QUAN_SIZE-1:0] = c2v_2[41];
assign v2c_2[41] = v2c_41_in2[QUAN_SIZE-1:0];
assign c2v_41_out3[QUAN_SIZE-1:0] = c2v_3[41];
assign v2c_3[41] = v2c_41_in3[QUAN_SIZE-1:0];
assign c2v_41_out4[QUAN_SIZE-1:0] = c2v_4[41];
assign v2c_4[41] = v2c_41_in4[QUAN_SIZE-1:0];
assign c2v_41_out5[QUAN_SIZE-1:0] = c2v_5[41];
assign v2c_5[41] = v2c_41_in5[QUAN_SIZE-1:0];
assign c2v_42_out0[QUAN_SIZE-1:0] = c2v_0[42];
assign v2c_0[42] = v2c_42_in0[QUAN_SIZE-1:0];
assign c2v_42_out1[QUAN_SIZE-1:0] = c2v_1[42];
assign v2c_1[42] = v2c_42_in1[QUAN_SIZE-1:0];
assign c2v_42_out2[QUAN_SIZE-1:0] = c2v_2[42];
assign v2c_2[42] = v2c_42_in2[QUAN_SIZE-1:0];
assign c2v_42_out3[QUAN_SIZE-1:0] = c2v_3[42];
assign v2c_3[42] = v2c_42_in3[QUAN_SIZE-1:0];
assign c2v_42_out4[QUAN_SIZE-1:0] = c2v_4[42];
assign v2c_4[42] = v2c_42_in4[QUAN_SIZE-1:0];
assign c2v_42_out5[QUAN_SIZE-1:0] = c2v_5[42];
assign v2c_5[42] = v2c_42_in5[QUAN_SIZE-1:0];
assign c2v_43_out0[QUAN_SIZE-1:0] = c2v_0[43];
assign v2c_0[43] = v2c_43_in0[QUAN_SIZE-1:0];
assign c2v_43_out1[QUAN_SIZE-1:0] = c2v_1[43];
assign v2c_1[43] = v2c_43_in1[QUAN_SIZE-1:0];
assign c2v_43_out2[QUAN_SIZE-1:0] = c2v_2[43];
assign v2c_2[43] = v2c_43_in2[QUAN_SIZE-1:0];
assign c2v_43_out3[QUAN_SIZE-1:0] = c2v_3[43];
assign v2c_3[43] = v2c_43_in3[QUAN_SIZE-1:0];
assign c2v_43_out4[QUAN_SIZE-1:0] = c2v_4[43];
assign v2c_4[43] = v2c_43_in4[QUAN_SIZE-1:0];
assign c2v_43_out5[QUAN_SIZE-1:0] = c2v_5[43];
assign v2c_5[43] = v2c_43_in5[QUAN_SIZE-1:0];
assign c2v_44_out0[QUAN_SIZE-1:0] = c2v_0[44];
assign v2c_0[44] = v2c_44_in0[QUAN_SIZE-1:0];
assign c2v_44_out1[QUAN_SIZE-1:0] = c2v_1[44];
assign v2c_1[44] = v2c_44_in1[QUAN_SIZE-1:0];
assign c2v_44_out2[QUAN_SIZE-1:0] = c2v_2[44];
assign v2c_2[44] = v2c_44_in2[QUAN_SIZE-1:0];
assign c2v_44_out3[QUAN_SIZE-1:0] = c2v_3[44];
assign v2c_3[44] = v2c_44_in3[QUAN_SIZE-1:0];
assign c2v_44_out4[QUAN_SIZE-1:0] = c2v_4[44];
assign v2c_4[44] = v2c_44_in4[QUAN_SIZE-1:0];
assign c2v_44_out5[QUAN_SIZE-1:0] = c2v_5[44];
assign v2c_5[44] = v2c_44_in5[QUAN_SIZE-1:0];
assign c2v_45_out0[QUAN_SIZE-1:0] = c2v_0[45];
assign v2c_0[45] = v2c_45_in0[QUAN_SIZE-1:0];
assign c2v_45_out1[QUAN_SIZE-1:0] = c2v_1[45];
assign v2c_1[45] = v2c_45_in1[QUAN_SIZE-1:0];
assign c2v_45_out2[QUAN_SIZE-1:0] = c2v_2[45];
assign v2c_2[45] = v2c_45_in2[QUAN_SIZE-1:0];
assign c2v_45_out3[QUAN_SIZE-1:0] = c2v_3[45];
assign v2c_3[45] = v2c_45_in3[QUAN_SIZE-1:0];
assign c2v_45_out4[QUAN_SIZE-1:0] = c2v_4[45];
assign v2c_4[45] = v2c_45_in4[QUAN_SIZE-1:0];
assign c2v_45_out5[QUAN_SIZE-1:0] = c2v_5[45];
assign v2c_5[45] = v2c_45_in5[QUAN_SIZE-1:0];
assign c2v_46_out0[QUAN_SIZE-1:0] = c2v_0[46];
assign v2c_0[46] = v2c_46_in0[QUAN_SIZE-1:0];
assign c2v_46_out1[QUAN_SIZE-1:0] = c2v_1[46];
assign v2c_1[46] = v2c_46_in1[QUAN_SIZE-1:0];
assign c2v_46_out2[QUAN_SIZE-1:0] = c2v_2[46];
assign v2c_2[46] = v2c_46_in2[QUAN_SIZE-1:0];
assign c2v_46_out3[QUAN_SIZE-1:0] = c2v_3[46];
assign v2c_3[46] = v2c_46_in3[QUAN_SIZE-1:0];
assign c2v_46_out4[QUAN_SIZE-1:0] = c2v_4[46];
assign v2c_4[46] = v2c_46_in4[QUAN_SIZE-1:0];
assign c2v_46_out5[QUAN_SIZE-1:0] = c2v_5[46];
assign v2c_5[46] = v2c_46_in5[QUAN_SIZE-1:0];
assign c2v_47_out0[QUAN_SIZE-1:0] = c2v_0[47];
assign v2c_0[47] = v2c_47_in0[QUAN_SIZE-1:0];
assign c2v_47_out1[QUAN_SIZE-1:0] = c2v_1[47];
assign v2c_1[47] = v2c_47_in1[QUAN_SIZE-1:0];
assign c2v_47_out2[QUAN_SIZE-1:0] = c2v_2[47];
assign v2c_2[47] = v2c_47_in2[QUAN_SIZE-1:0];
assign c2v_47_out3[QUAN_SIZE-1:0] = c2v_3[47];
assign v2c_3[47] = v2c_47_in3[QUAN_SIZE-1:0];
assign c2v_47_out4[QUAN_SIZE-1:0] = c2v_4[47];
assign v2c_4[47] = v2c_47_in4[QUAN_SIZE-1:0];
assign c2v_47_out5[QUAN_SIZE-1:0] = c2v_5[47];
assign v2c_5[47] = v2c_47_in5[QUAN_SIZE-1:0];
assign c2v_48_out0[QUAN_SIZE-1:0] = c2v_0[48];
assign v2c_0[48] = v2c_48_in0[QUAN_SIZE-1:0];
assign c2v_48_out1[QUAN_SIZE-1:0] = c2v_1[48];
assign v2c_1[48] = v2c_48_in1[QUAN_SIZE-1:0];
assign c2v_48_out2[QUAN_SIZE-1:0] = c2v_2[48];
assign v2c_2[48] = v2c_48_in2[QUAN_SIZE-1:0];
assign c2v_48_out3[QUAN_SIZE-1:0] = c2v_3[48];
assign v2c_3[48] = v2c_48_in3[QUAN_SIZE-1:0];
assign c2v_48_out4[QUAN_SIZE-1:0] = c2v_4[48];
assign v2c_4[48] = v2c_48_in4[QUAN_SIZE-1:0];
assign c2v_48_out5[QUAN_SIZE-1:0] = c2v_5[48];
assign v2c_5[48] = v2c_48_in5[QUAN_SIZE-1:0];
assign c2v_49_out0[QUAN_SIZE-1:0] = c2v_0[49];
assign v2c_0[49] = v2c_49_in0[QUAN_SIZE-1:0];
assign c2v_49_out1[QUAN_SIZE-1:0] = c2v_1[49];
assign v2c_1[49] = v2c_49_in1[QUAN_SIZE-1:0];
assign c2v_49_out2[QUAN_SIZE-1:0] = c2v_2[49];
assign v2c_2[49] = v2c_49_in2[QUAN_SIZE-1:0];
assign c2v_49_out3[QUAN_SIZE-1:0] = c2v_3[49];
assign v2c_3[49] = v2c_49_in3[QUAN_SIZE-1:0];
assign c2v_49_out4[QUAN_SIZE-1:0] = c2v_4[49];
assign v2c_4[49] = v2c_49_in4[QUAN_SIZE-1:0];
assign c2v_49_out5[QUAN_SIZE-1:0] = c2v_5[49];
assign v2c_5[49] = v2c_49_in5[QUAN_SIZE-1:0];
assign c2v_50_out0[QUAN_SIZE-1:0] = c2v_0[50];
assign v2c_0[50] = v2c_50_in0[QUAN_SIZE-1:0];
assign c2v_50_out1[QUAN_SIZE-1:0] = c2v_1[50];
assign v2c_1[50] = v2c_50_in1[QUAN_SIZE-1:0];
assign c2v_50_out2[QUAN_SIZE-1:0] = c2v_2[50];
assign v2c_2[50] = v2c_50_in2[QUAN_SIZE-1:0];
assign c2v_50_out3[QUAN_SIZE-1:0] = c2v_3[50];
assign v2c_3[50] = v2c_50_in3[QUAN_SIZE-1:0];
assign c2v_50_out4[QUAN_SIZE-1:0] = c2v_4[50];
assign v2c_4[50] = v2c_50_in4[QUAN_SIZE-1:0];
assign c2v_50_out5[QUAN_SIZE-1:0] = c2v_5[50];
assign v2c_5[50] = v2c_50_in5[QUAN_SIZE-1:0];
assign c2v_51_out0[QUAN_SIZE-1:0] = c2v_0[51];
assign v2c_0[51] = v2c_51_in0[QUAN_SIZE-1:0];
assign c2v_51_out1[QUAN_SIZE-1:0] = c2v_1[51];
assign v2c_1[51] = v2c_51_in1[QUAN_SIZE-1:0];
assign c2v_51_out2[QUAN_SIZE-1:0] = c2v_2[51];
assign v2c_2[51] = v2c_51_in2[QUAN_SIZE-1:0];
assign c2v_51_out3[QUAN_SIZE-1:0] = c2v_3[51];
assign v2c_3[51] = v2c_51_in3[QUAN_SIZE-1:0];
assign c2v_51_out4[QUAN_SIZE-1:0] = c2v_4[51];
assign v2c_4[51] = v2c_51_in4[QUAN_SIZE-1:0];
assign c2v_51_out5[QUAN_SIZE-1:0] = c2v_5[51];
assign v2c_5[51] = v2c_51_in5[QUAN_SIZE-1:0];
assign c2v_52_out0[QUAN_SIZE-1:0] = c2v_0[52];
assign v2c_0[52] = v2c_52_in0[QUAN_SIZE-1:0];
assign c2v_52_out1[QUAN_SIZE-1:0] = c2v_1[52];
assign v2c_1[52] = v2c_52_in1[QUAN_SIZE-1:0];
assign c2v_52_out2[QUAN_SIZE-1:0] = c2v_2[52];
assign v2c_2[52] = v2c_52_in2[QUAN_SIZE-1:0];
assign c2v_52_out3[QUAN_SIZE-1:0] = c2v_3[52];
assign v2c_3[52] = v2c_52_in3[QUAN_SIZE-1:0];
assign c2v_52_out4[QUAN_SIZE-1:0] = c2v_4[52];
assign v2c_4[52] = v2c_52_in4[QUAN_SIZE-1:0];
assign c2v_52_out5[QUAN_SIZE-1:0] = c2v_5[52];
assign v2c_5[52] = v2c_52_in5[QUAN_SIZE-1:0];
assign c2v_53_out0[QUAN_SIZE-1:0] = c2v_0[53];
assign v2c_0[53] = v2c_53_in0[QUAN_SIZE-1:0];
assign c2v_53_out1[QUAN_SIZE-1:0] = c2v_1[53];
assign v2c_1[53] = v2c_53_in1[QUAN_SIZE-1:0];
assign c2v_53_out2[QUAN_SIZE-1:0] = c2v_2[53];
assign v2c_2[53] = v2c_53_in2[QUAN_SIZE-1:0];
assign c2v_53_out3[QUAN_SIZE-1:0] = c2v_3[53];
assign v2c_3[53] = v2c_53_in3[QUAN_SIZE-1:0];
assign c2v_53_out4[QUAN_SIZE-1:0] = c2v_4[53];
assign v2c_4[53] = v2c_53_in4[QUAN_SIZE-1:0];
assign c2v_53_out5[QUAN_SIZE-1:0] = c2v_5[53];
assign v2c_5[53] = v2c_53_in5[QUAN_SIZE-1:0];
assign c2v_54_out0[QUAN_SIZE-1:0] = c2v_0[54];
assign v2c_0[54] = v2c_54_in0[QUAN_SIZE-1:0];
assign c2v_54_out1[QUAN_SIZE-1:0] = c2v_1[54];
assign v2c_1[54] = v2c_54_in1[QUAN_SIZE-1:0];
assign c2v_54_out2[QUAN_SIZE-1:0] = c2v_2[54];
assign v2c_2[54] = v2c_54_in2[QUAN_SIZE-1:0];
assign c2v_54_out3[QUAN_SIZE-1:0] = c2v_3[54];
assign v2c_3[54] = v2c_54_in3[QUAN_SIZE-1:0];
assign c2v_54_out4[QUAN_SIZE-1:0] = c2v_4[54];
assign v2c_4[54] = v2c_54_in4[QUAN_SIZE-1:0];
assign c2v_54_out5[QUAN_SIZE-1:0] = c2v_5[54];
assign v2c_5[54] = v2c_54_in5[QUAN_SIZE-1:0];
assign c2v_55_out0[QUAN_SIZE-1:0] = c2v_0[55];
assign v2c_0[55] = v2c_55_in0[QUAN_SIZE-1:0];
assign c2v_55_out1[QUAN_SIZE-1:0] = c2v_1[55];
assign v2c_1[55] = v2c_55_in1[QUAN_SIZE-1:0];
assign c2v_55_out2[QUAN_SIZE-1:0] = c2v_2[55];
assign v2c_2[55] = v2c_55_in2[QUAN_SIZE-1:0];
assign c2v_55_out3[QUAN_SIZE-1:0] = c2v_3[55];
assign v2c_3[55] = v2c_55_in3[QUAN_SIZE-1:0];
assign c2v_55_out4[QUAN_SIZE-1:0] = c2v_4[55];
assign v2c_4[55] = v2c_55_in4[QUAN_SIZE-1:0];
assign c2v_55_out5[QUAN_SIZE-1:0] = c2v_5[55];
assign v2c_5[55] = v2c_55_in5[QUAN_SIZE-1:0];
assign c2v_56_out0[QUAN_SIZE-1:0] = c2v_0[56];
assign v2c_0[56] = v2c_56_in0[QUAN_SIZE-1:0];
assign c2v_56_out1[QUAN_SIZE-1:0] = c2v_1[56];
assign v2c_1[56] = v2c_56_in1[QUAN_SIZE-1:0];
assign c2v_56_out2[QUAN_SIZE-1:0] = c2v_2[56];
assign v2c_2[56] = v2c_56_in2[QUAN_SIZE-1:0];
assign c2v_56_out3[QUAN_SIZE-1:0] = c2v_3[56];
assign v2c_3[56] = v2c_56_in3[QUAN_SIZE-1:0];
assign c2v_56_out4[QUAN_SIZE-1:0] = c2v_4[56];
assign v2c_4[56] = v2c_56_in4[QUAN_SIZE-1:0];
assign c2v_56_out5[QUAN_SIZE-1:0] = c2v_5[56];
assign v2c_5[56] = v2c_56_in5[QUAN_SIZE-1:0];
assign c2v_57_out0[QUAN_SIZE-1:0] = c2v_0[57];
assign v2c_0[57] = v2c_57_in0[QUAN_SIZE-1:0];
assign c2v_57_out1[QUAN_SIZE-1:0] = c2v_1[57];
assign v2c_1[57] = v2c_57_in1[QUAN_SIZE-1:0];
assign c2v_57_out2[QUAN_SIZE-1:0] = c2v_2[57];
assign v2c_2[57] = v2c_57_in2[QUAN_SIZE-1:0];
assign c2v_57_out3[QUAN_SIZE-1:0] = c2v_3[57];
assign v2c_3[57] = v2c_57_in3[QUAN_SIZE-1:0];
assign c2v_57_out4[QUAN_SIZE-1:0] = c2v_4[57];
assign v2c_4[57] = v2c_57_in4[QUAN_SIZE-1:0];
assign c2v_57_out5[QUAN_SIZE-1:0] = c2v_5[57];
assign v2c_5[57] = v2c_57_in5[QUAN_SIZE-1:0];
assign c2v_58_out0[QUAN_SIZE-1:0] = c2v_0[58];
assign v2c_0[58] = v2c_58_in0[QUAN_SIZE-1:0];
assign c2v_58_out1[QUAN_SIZE-1:0] = c2v_1[58];
assign v2c_1[58] = v2c_58_in1[QUAN_SIZE-1:0];
assign c2v_58_out2[QUAN_SIZE-1:0] = c2v_2[58];
assign v2c_2[58] = v2c_58_in2[QUAN_SIZE-1:0];
assign c2v_58_out3[QUAN_SIZE-1:0] = c2v_3[58];
assign v2c_3[58] = v2c_58_in3[QUAN_SIZE-1:0];
assign c2v_58_out4[QUAN_SIZE-1:0] = c2v_4[58];
assign v2c_4[58] = v2c_58_in4[QUAN_SIZE-1:0];
assign c2v_58_out5[QUAN_SIZE-1:0] = c2v_5[58];
assign v2c_5[58] = v2c_58_in5[QUAN_SIZE-1:0];
assign c2v_59_out0[QUAN_SIZE-1:0] = c2v_0[59];
assign v2c_0[59] = v2c_59_in0[QUAN_SIZE-1:0];
assign c2v_59_out1[QUAN_SIZE-1:0] = c2v_1[59];
assign v2c_1[59] = v2c_59_in1[QUAN_SIZE-1:0];
assign c2v_59_out2[QUAN_SIZE-1:0] = c2v_2[59];
assign v2c_2[59] = v2c_59_in2[QUAN_SIZE-1:0];
assign c2v_59_out3[QUAN_SIZE-1:0] = c2v_3[59];
assign v2c_3[59] = v2c_59_in3[QUAN_SIZE-1:0];
assign c2v_59_out4[QUAN_SIZE-1:0] = c2v_4[59];
assign v2c_4[59] = v2c_59_in4[QUAN_SIZE-1:0];
assign c2v_59_out5[QUAN_SIZE-1:0] = c2v_5[59];
assign v2c_5[59] = v2c_59_in5[QUAN_SIZE-1:0];
assign c2v_60_out0[QUAN_SIZE-1:0] = c2v_0[60];
assign v2c_0[60] = v2c_60_in0[QUAN_SIZE-1:0];
assign c2v_60_out1[QUAN_SIZE-1:0] = c2v_1[60];
assign v2c_1[60] = v2c_60_in1[QUAN_SIZE-1:0];
assign c2v_60_out2[QUAN_SIZE-1:0] = c2v_2[60];
assign v2c_2[60] = v2c_60_in2[QUAN_SIZE-1:0];
assign c2v_60_out3[QUAN_SIZE-1:0] = c2v_3[60];
assign v2c_3[60] = v2c_60_in3[QUAN_SIZE-1:0];
assign c2v_60_out4[QUAN_SIZE-1:0] = c2v_4[60];
assign v2c_4[60] = v2c_60_in4[QUAN_SIZE-1:0];
assign c2v_60_out5[QUAN_SIZE-1:0] = c2v_5[60];
assign v2c_5[60] = v2c_60_in5[QUAN_SIZE-1:0];
assign c2v_61_out0[QUAN_SIZE-1:0] = c2v_0[61];
assign v2c_0[61] = v2c_61_in0[QUAN_SIZE-1:0];
assign c2v_61_out1[QUAN_SIZE-1:0] = c2v_1[61];
assign v2c_1[61] = v2c_61_in1[QUAN_SIZE-1:0];
assign c2v_61_out2[QUAN_SIZE-1:0] = c2v_2[61];
assign v2c_2[61] = v2c_61_in2[QUAN_SIZE-1:0];
assign c2v_61_out3[QUAN_SIZE-1:0] = c2v_3[61];
assign v2c_3[61] = v2c_61_in3[QUAN_SIZE-1:0];
assign c2v_61_out4[QUAN_SIZE-1:0] = c2v_4[61];
assign v2c_4[61] = v2c_61_in4[QUAN_SIZE-1:0];
assign c2v_61_out5[QUAN_SIZE-1:0] = c2v_5[61];
assign v2c_5[61] = v2c_61_in5[QUAN_SIZE-1:0];
assign c2v_62_out0[QUAN_SIZE-1:0] = c2v_0[62];
assign v2c_0[62] = v2c_62_in0[QUAN_SIZE-1:0];
assign c2v_62_out1[QUAN_SIZE-1:0] = c2v_1[62];
assign v2c_1[62] = v2c_62_in1[QUAN_SIZE-1:0];
assign c2v_62_out2[QUAN_SIZE-1:0] = c2v_2[62];
assign v2c_2[62] = v2c_62_in2[QUAN_SIZE-1:0];
assign c2v_62_out3[QUAN_SIZE-1:0] = c2v_3[62];
assign v2c_3[62] = v2c_62_in3[QUAN_SIZE-1:0];
assign c2v_62_out4[QUAN_SIZE-1:0] = c2v_4[62];
assign v2c_4[62] = v2c_62_in4[QUAN_SIZE-1:0];
assign c2v_62_out5[QUAN_SIZE-1:0] = c2v_5[62];
assign v2c_5[62] = v2c_62_in5[QUAN_SIZE-1:0];
assign c2v_63_out0[QUAN_SIZE-1:0] = c2v_0[63];
assign v2c_0[63] = v2c_63_in0[QUAN_SIZE-1:0];
assign c2v_63_out1[QUAN_SIZE-1:0] = c2v_1[63];
assign v2c_1[63] = v2c_63_in1[QUAN_SIZE-1:0];
assign c2v_63_out2[QUAN_SIZE-1:0] = c2v_2[63];
assign v2c_2[63] = v2c_63_in2[QUAN_SIZE-1:0];
assign c2v_63_out3[QUAN_SIZE-1:0] = c2v_3[63];
assign v2c_3[63] = v2c_63_in3[QUAN_SIZE-1:0];
assign c2v_63_out4[QUAN_SIZE-1:0] = c2v_4[63];
assign v2c_4[63] = v2c_63_in4[QUAN_SIZE-1:0];
assign c2v_63_out5[QUAN_SIZE-1:0] = c2v_5[63];
assign v2c_5[63] = v2c_63_in5[QUAN_SIZE-1:0];
assign c2v_64_out0[QUAN_SIZE-1:0] = c2v_0[64];
assign v2c_0[64] = v2c_64_in0[QUAN_SIZE-1:0];
assign c2v_64_out1[QUAN_SIZE-1:0] = c2v_1[64];
assign v2c_1[64] = v2c_64_in1[QUAN_SIZE-1:0];
assign c2v_64_out2[QUAN_SIZE-1:0] = c2v_2[64];
assign v2c_2[64] = v2c_64_in2[QUAN_SIZE-1:0];
assign c2v_64_out3[QUAN_SIZE-1:0] = c2v_3[64];
assign v2c_3[64] = v2c_64_in3[QUAN_SIZE-1:0];
assign c2v_64_out4[QUAN_SIZE-1:0] = c2v_4[64];
assign v2c_4[64] = v2c_64_in4[QUAN_SIZE-1:0];
assign c2v_64_out5[QUAN_SIZE-1:0] = c2v_5[64];
assign v2c_5[64] = v2c_64_in5[QUAN_SIZE-1:0];
assign c2v_65_out0[QUAN_SIZE-1:0] = c2v_0[65];
assign v2c_0[65] = v2c_65_in0[QUAN_SIZE-1:0];
assign c2v_65_out1[QUAN_SIZE-1:0] = c2v_1[65];
assign v2c_1[65] = v2c_65_in1[QUAN_SIZE-1:0];
assign c2v_65_out2[QUAN_SIZE-1:0] = c2v_2[65];
assign v2c_2[65] = v2c_65_in2[QUAN_SIZE-1:0];
assign c2v_65_out3[QUAN_SIZE-1:0] = c2v_3[65];
assign v2c_3[65] = v2c_65_in3[QUAN_SIZE-1:0];
assign c2v_65_out4[QUAN_SIZE-1:0] = c2v_4[65];
assign v2c_4[65] = v2c_65_in4[QUAN_SIZE-1:0];
assign c2v_65_out5[QUAN_SIZE-1:0] = c2v_5[65];
assign v2c_5[65] = v2c_65_in5[QUAN_SIZE-1:0];
assign c2v_66_out0[QUAN_SIZE-1:0] = c2v_0[66];
assign v2c_0[66] = v2c_66_in0[QUAN_SIZE-1:0];
assign c2v_66_out1[QUAN_SIZE-1:0] = c2v_1[66];
assign v2c_1[66] = v2c_66_in1[QUAN_SIZE-1:0];
assign c2v_66_out2[QUAN_SIZE-1:0] = c2v_2[66];
assign v2c_2[66] = v2c_66_in2[QUAN_SIZE-1:0];
assign c2v_66_out3[QUAN_SIZE-1:0] = c2v_3[66];
assign v2c_3[66] = v2c_66_in3[QUAN_SIZE-1:0];
assign c2v_66_out4[QUAN_SIZE-1:0] = c2v_4[66];
assign v2c_4[66] = v2c_66_in4[QUAN_SIZE-1:0];
assign c2v_66_out5[QUAN_SIZE-1:0] = c2v_5[66];
assign v2c_5[66] = v2c_66_in5[QUAN_SIZE-1:0];
assign c2v_67_out0[QUAN_SIZE-1:0] = c2v_0[67];
assign v2c_0[67] = v2c_67_in0[QUAN_SIZE-1:0];
assign c2v_67_out1[QUAN_SIZE-1:0] = c2v_1[67];
assign v2c_1[67] = v2c_67_in1[QUAN_SIZE-1:0];
assign c2v_67_out2[QUAN_SIZE-1:0] = c2v_2[67];
assign v2c_2[67] = v2c_67_in2[QUAN_SIZE-1:0];
assign c2v_67_out3[QUAN_SIZE-1:0] = c2v_3[67];
assign v2c_3[67] = v2c_67_in3[QUAN_SIZE-1:0];
assign c2v_67_out4[QUAN_SIZE-1:0] = c2v_4[67];
assign v2c_4[67] = v2c_67_in4[QUAN_SIZE-1:0];
assign c2v_67_out5[QUAN_SIZE-1:0] = c2v_5[67];
assign v2c_5[67] = v2c_67_in5[QUAN_SIZE-1:0];
assign c2v_68_out0[QUAN_SIZE-1:0] = c2v_0[68];
assign v2c_0[68] = v2c_68_in0[QUAN_SIZE-1:0];
assign c2v_68_out1[QUAN_SIZE-1:0] = c2v_1[68];
assign v2c_1[68] = v2c_68_in1[QUAN_SIZE-1:0];
assign c2v_68_out2[QUAN_SIZE-1:0] = c2v_2[68];
assign v2c_2[68] = v2c_68_in2[QUAN_SIZE-1:0];
assign c2v_68_out3[QUAN_SIZE-1:0] = c2v_3[68];
assign v2c_3[68] = v2c_68_in3[QUAN_SIZE-1:0];
assign c2v_68_out4[QUAN_SIZE-1:0] = c2v_4[68];
assign v2c_4[68] = v2c_68_in4[QUAN_SIZE-1:0];
assign c2v_68_out5[QUAN_SIZE-1:0] = c2v_5[68];
assign v2c_5[68] = v2c_68_in5[QUAN_SIZE-1:0];
assign c2v_69_out0[QUAN_SIZE-1:0] = c2v_0[69];
assign v2c_0[69] = v2c_69_in0[QUAN_SIZE-1:0];
assign c2v_69_out1[QUAN_SIZE-1:0] = c2v_1[69];
assign v2c_1[69] = v2c_69_in1[QUAN_SIZE-1:0];
assign c2v_69_out2[QUAN_SIZE-1:0] = c2v_2[69];
assign v2c_2[69] = v2c_69_in2[QUAN_SIZE-1:0];
assign c2v_69_out3[QUAN_SIZE-1:0] = c2v_3[69];
assign v2c_3[69] = v2c_69_in3[QUAN_SIZE-1:0];
assign c2v_69_out4[QUAN_SIZE-1:0] = c2v_4[69];
assign v2c_4[69] = v2c_69_in4[QUAN_SIZE-1:0];
assign c2v_69_out5[QUAN_SIZE-1:0] = c2v_5[69];
assign v2c_5[69] = v2c_69_in5[QUAN_SIZE-1:0];
assign c2v_70_out0[QUAN_SIZE-1:0] = c2v_0[70];
assign v2c_0[70] = v2c_70_in0[QUAN_SIZE-1:0];
assign c2v_70_out1[QUAN_SIZE-1:0] = c2v_1[70];
assign v2c_1[70] = v2c_70_in1[QUAN_SIZE-1:0];
assign c2v_70_out2[QUAN_SIZE-1:0] = c2v_2[70];
assign v2c_2[70] = v2c_70_in2[QUAN_SIZE-1:0];
assign c2v_70_out3[QUAN_SIZE-1:0] = c2v_3[70];
assign v2c_3[70] = v2c_70_in3[QUAN_SIZE-1:0];
assign c2v_70_out4[QUAN_SIZE-1:0] = c2v_4[70];
assign v2c_4[70] = v2c_70_in4[QUAN_SIZE-1:0];
assign c2v_70_out5[QUAN_SIZE-1:0] = c2v_5[70];
assign v2c_5[70] = v2c_70_in5[QUAN_SIZE-1:0];
assign c2v_71_out0[QUAN_SIZE-1:0] = c2v_0[71];
assign v2c_0[71] = v2c_71_in0[QUAN_SIZE-1:0];
assign c2v_71_out1[QUAN_SIZE-1:0] = c2v_1[71];
assign v2c_1[71] = v2c_71_in1[QUAN_SIZE-1:0];
assign c2v_71_out2[QUAN_SIZE-1:0] = c2v_2[71];
assign v2c_2[71] = v2c_71_in2[QUAN_SIZE-1:0];
assign c2v_71_out3[QUAN_SIZE-1:0] = c2v_3[71];
assign v2c_3[71] = v2c_71_in3[QUAN_SIZE-1:0];
assign c2v_71_out4[QUAN_SIZE-1:0] = c2v_4[71];
assign v2c_4[71] = v2c_71_in4[QUAN_SIZE-1:0];
assign c2v_71_out5[QUAN_SIZE-1:0] = c2v_5[71];
assign v2c_5[71] = v2c_71_in5[QUAN_SIZE-1:0];
assign c2v_72_out0[QUAN_SIZE-1:0] = c2v_0[72];
assign v2c_0[72] = v2c_72_in0[QUAN_SIZE-1:0];
assign c2v_72_out1[QUAN_SIZE-1:0] = c2v_1[72];
assign v2c_1[72] = v2c_72_in1[QUAN_SIZE-1:0];
assign c2v_72_out2[QUAN_SIZE-1:0] = c2v_2[72];
assign v2c_2[72] = v2c_72_in2[QUAN_SIZE-1:0];
assign c2v_72_out3[QUAN_SIZE-1:0] = c2v_3[72];
assign v2c_3[72] = v2c_72_in3[QUAN_SIZE-1:0];
assign c2v_72_out4[QUAN_SIZE-1:0] = c2v_4[72];
assign v2c_4[72] = v2c_72_in4[QUAN_SIZE-1:0];
assign c2v_72_out5[QUAN_SIZE-1:0] = c2v_5[72];
assign v2c_5[72] = v2c_72_in5[QUAN_SIZE-1:0];
assign c2v_73_out0[QUAN_SIZE-1:0] = c2v_0[73];
assign v2c_0[73] = v2c_73_in0[QUAN_SIZE-1:0];
assign c2v_73_out1[QUAN_SIZE-1:0] = c2v_1[73];
assign v2c_1[73] = v2c_73_in1[QUAN_SIZE-1:0];
assign c2v_73_out2[QUAN_SIZE-1:0] = c2v_2[73];
assign v2c_2[73] = v2c_73_in2[QUAN_SIZE-1:0];
assign c2v_73_out3[QUAN_SIZE-1:0] = c2v_3[73];
assign v2c_3[73] = v2c_73_in3[QUAN_SIZE-1:0];
assign c2v_73_out4[QUAN_SIZE-1:0] = c2v_4[73];
assign v2c_4[73] = v2c_73_in4[QUAN_SIZE-1:0];
assign c2v_73_out5[QUAN_SIZE-1:0] = c2v_5[73];
assign v2c_5[73] = v2c_73_in5[QUAN_SIZE-1:0];
assign c2v_74_out0[QUAN_SIZE-1:0] = c2v_0[74];
assign v2c_0[74] = v2c_74_in0[QUAN_SIZE-1:0];
assign c2v_74_out1[QUAN_SIZE-1:0] = c2v_1[74];
assign v2c_1[74] = v2c_74_in1[QUAN_SIZE-1:0];
assign c2v_74_out2[QUAN_SIZE-1:0] = c2v_2[74];
assign v2c_2[74] = v2c_74_in2[QUAN_SIZE-1:0];
assign c2v_74_out3[QUAN_SIZE-1:0] = c2v_3[74];
assign v2c_3[74] = v2c_74_in3[QUAN_SIZE-1:0];
assign c2v_74_out4[QUAN_SIZE-1:0] = c2v_4[74];
assign v2c_4[74] = v2c_74_in4[QUAN_SIZE-1:0];
assign c2v_74_out5[QUAN_SIZE-1:0] = c2v_5[74];
assign v2c_5[74] = v2c_74_in5[QUAN_SIZE-1:0];
assign c2v_75_out0[QUAN_SIZE-1:0] = c2v_0[75];
assign v2c_0[75] = v2c_75_in0[QUAN_SIZE-1:0];
assign c2v_75_out1[QUAN_SIZE-1:0] = c2v_1[75];
assign v2c_1[75] = v2c_75_in1[QUAN_SIZE-1:0];
assign c2v_75_out2[QUAN_SIZE-1:0] = c2v_2[75];
assign v2c_2[75] = v2c_75_in2[QUAN_SIZE-1:0];
assign c2v_75_out3[QUAN_SIZE-1:0] = c2v_3[75];
assign v2c_3[75] = v2c_75_in3[QUAN_SIZE-1:0];
assign c2v_75_out4[QUAN_SIZE-1:0] = c2v_4[75];
assign v2c_4[75] = v2c_75_in4[QUAN_SIZE-1:0];
assign c2v_75_out5[QUAN_SIZE-1:0] = c2v_5[75];
assign v2c_5[75] = v2c_75_in5[QUAN_SIZE-1:0];
assign c2v_76_out0[QUAN_SIZE-1:0] = c2v_0[76];
assign v2c_0[76] = v2c_76_in0[QUAN_SIZE-1:0];
assign c2v_76_out1[QUAN_SIZE-1:0] = c2v_1[76];
assign v2c_1[76] = v2c_76_in1[QUAN_SIZE-1:0];
assign c2v_76_out2[QUAN_SIZE-1:0] = c2v_2[76];
assign v2c_2[76] = v2c_76_in2[QUAN_SIZE-1:0];
assign c2v_76_out3[QUAN_SIZE-1:0] = c2v_3[76];
assign v2c_3[76] = v2c_76_in3[QUAN_SIZE-1:0];
assign c2v_76_out4[QUAN_SIZE-1:0] = c2v_4[76];
assign v2c_4[76] = v2c_76_in4[QUAN_SIZE-1:0];
assign c2v_76_out5[QUAN_SIZE-1:0] = c2v_5[76];
assign v2c_5[76] = v2c_76_in5[QUAN_SIZE-1:0];
assign c2v_77_out0[QUAN_SIZE-1:0] = c2v_0[77];
assign v2c_0[77] = v2c_77_in0[QUAN_SIZE-1:0];
assign c2v_77_out1[QUAN_SIZE-1:0] = c2v_1[77];
assign v2c_1[77] = v2c_77_in1[QUAN_SIZE-1:0];
assign c2v_77_out2[QUAN_SIZE-1:0] = c2v_2[77];
assign v2c_2[77] = v2c_77_in2[QUAN_SIZE-1:0];
assign c2v_77_out3[QUAN_SIZE-1:0] = c2v_3[77];
assign v2c_3[77] = v2c_77_in3[QUAN_SIZE-1:0];
assign c2v_77_out4[QUAN_SIZE-1:0] = c2v_4[77];
assign v2c_4[77] = v2c_77_in4[QUAN_SIZE-1:0];
assign c2v_77_out5[QUAN_SIZE-1:0] = c2v_5[77];
assign v2c_5[77] = v2c_77_in5[QUAN_SIZE-1:0];
assign c2v_78_out0[QUAN_SIZE-1:0] = c2v_0[78];
assign v2c_0[78] = v2c_78_in0[QUAN_SIZE-1:0];
assign c2v_78_out1[QUAN_SIZE-1:0] = c2v_1[78];
assign v2c_1[78] = v2c_78_in1[QUAN_SIZE-1:0];
assign c2v_78_out2[QUAN_SIZE-1:0] = c2v_2[78];
assign v2c_2[78] = v2c_78_in2[QUAN_SIZE-1:0];
assign c2v_78_out3[QUAN_SIZE-1:0] = c2v_3[78];
assign v2c_3[78] = v2c_78_in3[QUAN_SIZE-1:0];
assign c2v_78_out4[QUAN_SIZE-1:0] = c2v_4[78];
assign v2c_4[78] = v2c_78_in4[QUAN_SIZE-1:0];
assign c2v_78_out5[QUAN_SIZE-1:0] = c2v_5[78];
assign v2c_5[78] = v2c_78_in5[QUAN_SIZE-1:0];
assign c2v_79_out0[QUAN_SIZE-1:0] = c2v_0[79];
assign v2c_0[79] = v2c_79_in0[QUAN_SIZE-1:0];
assign c2v_79_out1[QUAN_SIZE-1:0] = c2v_1[79];
assign v2c_1[79] = v2c_79_in1[QUAN_SIZE-1:0];
assign c2v_79_out2[QUAN_SIZE-1:0] = c2v_2[79];
assign v2c_2[79] = v2c_79_in2[QUAN_SIZE-1:0];
assign c2v_79_out3[QUAN_SIZE-1:0] = c2v_3[79];
assign v2c_3[79] = v2c_79_in3[QUAN_SIZE-1:0];
assign c2v_79_out4[QUAN_SIZE-1:0] = c2v_4[79];
assign v2c_4[79] = v2c_79_in4[QUAN_SIZE-1:0];
assign c2v_79_out5[QUAN_SIZE-1:0] = c2v_5[79];
assign v2c_5[79] = v2c_79_in5[QUAN_SIZE-1:0];
assign c2v_80_out0[QUAN_SIZE-1:0] = c2v_0[80];
assign v2c_0[80] = v2c_80_in0[QUAN_SIZE-1:0];
assign c2v_80_out1[QUAN_SIZE-1:0] = c2v_1[80];
assign v2c_1[80] = v2c_80_in1[QUAN_SIZE-1:0];
assign c2v_80_out2[QUAN_SIZE-1:0] = c2v_2[80];
assign v2c_2[80] = v2c_80_in2[QUAN_SIZE-1:0];
assign c2v_80_out3[QUAN_SIZE-1:0] = c2v_3[80];
assign v2c_3[80] = v2c_80_in3[QUAN_SIZE-1:0];
assign c2v_80_out4[QUAN_SIZE-1:0] = c2v_4[80];
assign v2c_4[80] = v2c_80_in4[QUAN_SIZE-1:0];
assign c2v_80_out5[QUAN_SIZE-1:0] = c2v_5[80];
assign v2c_5[80] = v2c_80_in5[QUAN_SIZE-1:0];
assign c2v_81_out0[QUAN_SIZE-1:0] = c2v_0[81];
assign v2c_0[81] = v2c_81_in0[QUAN_SIZE-1:0];
assign c2v_81_out1[QUAN_SIZE-1:0] = c2v_1[81];
assign v2c_1[81] = v2c_81_in1[QUAN_SIZE-1:0];
assign c2v_81_out2[QUAN_SIZE-1:0] = c2v_2[81];
assign v2c_2[81] = v2c_81_in2[QUAN_SIZE-1:0];
assign c2v_81_out3[QUAN_SIZE-1:0] = c2v_3[81];
assign v2c_3[81] = v2c_81_in3[QUAN_SIZE-1:0];
assign c2v_81_out4[QUAN_SIZE-1:0] = c2v_4[81];
assign v2c_4[81] = v2c_81_in4[QUAN_SIZE-1:0];
assign c2v_81_out5[QUAN_SIZE-1:0] = c2v_5[81];
assign v2c_5[81] = v2c_81_in5[QUAN_SIZE-1:0];
assign c2v_82_out0[QUAN_SIZE-1:0] = c2v_0[82];
assign v2c_0[82] = v2c_82_in0[QUAN_SIZE-1:0];
assign c2v_82_out1[QUAN_SIZE-1:0] = c2v_1[82];
assign v2c_1[82] = v2c_82_in1[QUAN_SIZE-1:0];
assign c2v_82_out2[QUAN_SIZE-1:0] = c2v_2[82];
assign v2c_2[82] = v2c_82_in2[QUAN_SIZE-1:0];
assign c2v_82_out3[QUAN_SIZE-1:0] = c2v_3[82];
assign v2c_3[82] = v2c_82_in3[QUAN_SIZE-1:0];
assign c2v_82_out4[QUAN_SIZE-1:0] = c2v_4[82];
assign v2c_4[82] = v2c_82_in4[QUAN_SIZE-1:0];
assign c2v_82_out5[QUAN_SIZE-1:0] = c2v_5[82];
assign v2c_5[82] = v2c_82_in5[QUAN_SIZE-1:0];
assign c2v_83_out0[QUAN_SIZE-1:0] = c2v_0[83];
assign v2c_0[83] = v2c_83_in0[QUAN_SIZE-1:0];
assign c2v_83_out1[QUAN_SIZE-1:0] = c2v_1[83];
assign v2c_1[83] = v2c_83_in1[QUAN_SIZE-1:0];
assign c2v_83_out2[QUAN_SIZE-1:0] = c2v_2[83];
assign v2c_2[83] = v2c_83_in2[QUAN_SIZE-1:0];
assign c2v_83_out3[QUAN_SIZE-1:0] = c2v_3[83];
assign v2c_3[83] = v2c_83_in3[QUAN_SIZE-1:0];
assign c2v_83_out4[QUAN_SIZE-1:0] = c2v_4[83];
assign v2c_4[83] = v2c_83_in4[QUAN_SIZE-1:0];
assign c2v_83_out5[QUAN_SIZE-1:0] = c2v_5[83];
assign v2c_5[83] = v2c_83_in5[QUAN_SIZE-1:0];
assign c2v_84_out0[QUAN_SIZE-1:0] = c2v_0[84];
assign v2c_0[84] = v2c_84_in0[QUAN_SIZE-1:0];
assign c2v_84_out1[QUAN_SIZE-1:0] = c2v_1[84];
assign v2c_1[84] = v2c_84_in1[QUAN_SIZE-1:0];
assign c2v_84_out2[QUAN_SIZE-1:0] = c2v_2[84];
assign v2c_2[84] = v2c_84_in2[QUAN_SIZE-1:0];
assign c2v_84_out3[QUAN_SIZE-1:0] = c2v_3[84];
assign v2c_3[84] = v2c_84_in3[QUAN_SIZE-1:0];
assign c2v_84_out4[QUAN_SIZE-1:0] = c2v_4[84];
assign v2c_4[84] = v2c_84_in4[QUAN_SIZE-1:0];
assign c2v_84_out5[QUAN_SIZE-1:0] = c2v_5[84];
assign v2c_5[84] = v2c_84_in5[QUAN_SIZE-1:0];
assign c2v_85_out0[QUAN_SIZE-1:0] = c2v_0[85];
assign v2c_0[85] = v2c_85_in0[QUAN_SIZE-1:0];
assign c2v_85_out1[QUAN_SIZE-1:0] = c2v_1[85];
assign v2c_1[85] = v2c_85_in1[QUAN_SIZE-1:0];
assign c2v_85_out2[QUAN_SIZE-1:0] = c2v_2[85];
assign v2c_2[85] = v2c_85_in2[QUAN_SIZE-1:0];
assign c2v_85_out3[QUAN_SIZE-1:0] = c2v_3[85];
assign v2c_3[85] = v2c_85_in3[QUAN_SIZE-1:0];
assign c2v_85_out4[QUAN_SIZE-1:0] = c2v_4[85];
assign v2c_4[85] = v2c_85_in4[QUAN_SIZE-1:0];
assign c2v_85_out5[QUAN_SIZE-1:0] = c2v_5[85];
assign v2c_5[85] = v2c_85_in5[QUAN_SIZE-1:0];
assign c2v_86_out0[QUAN_SIZE-1:0] = c2v_0[86];
assign v2c_0[86] = v2c_86_in0[QUAN_SIZE-1:0];
assign c2v_86_out1[QUAN_SIZE-1:0] = c2v_1[86];
assign v2c_1[86] = v2c_86_in1[QUAN_SIZE-1:0];
assign c2v_86_out2[QUAN_SIZE-1:0] = c2v_2[86];
assign v2c_2[86] = v2c_86_in2[QUAN_SIZE-1:0];
assign c2v_86_out3[QUAN_SIZE-1:0] = c2v_3[86];
assign v2c_3[86] = v2c_86_in3[QUAN_SIZE-1:0];
assign c2v_86_out4[QUAN_SIZE-1:0] = c2v_4[86];
assign v2c_4[86] = v2c_86_in4[QUAN_SIZE-1:0];
assign c2v_86_out5[QUAN_SIZE-1:0] = c2v_5[86];
assign v2c_5[86] = v2c_86_in5[QUAN_SIZE-1:0];
assign c2v_87_out0[QUAN_SIZE-1:0] = c2v_0[87];
assign v2c_0[87] = v2c_87_in0[QUAN_SIZE-1:0];
assign c2v_87_out1[QUAN_SIZE-1:0] = c2v_1[87];
assign v2c_1[87] = v2c_87_in1[QUAN_SIZE-1:0];
assign c2v_87_out2[QUAN_SIZE-1:0] = c2v_2[87];
assign v2c_2[87] = v2c_87_in2[QUAN_SIZE-1:0];
assign c2v_87_out3[QUAN_SIZE-1:0] = c2v_3[87];
assign v2c_3[87] = v2c_87_in3[QUAN_SIZE-1:0];
assign c2v_87_out4[QUAN_SIZE-1:0] = c2v_4[87];
assign v2c_4[87] = v2c_87_in4[QUAN_SIZE-1:0];
assign c2v_87_out5[QUAN_SIZE-1:0] = c2v_5[87];
assign v2c_5[87] = v2c_87_in5[QUAN_SIZE-1:0];
assign c2v_88_out0[QUAN_SIZE-1:0] = c2v_0[88];
assign v2c_0[88] = v2c_88_in0[QUAN_SIZE-1:0];
assign c2v_88_out1[QUAN_SIZE-1:0] = c2v_1[88];
assign v2c_1[88] = v2c_88_in1[QUAN_SIZE-1:0];
assign c2v_88_out2[QUAN_SIZE-1:0] = c2v_2[88];
assign v2c_2[88] = v2c_88_in2[QUAN_SIZE-1:0];
assign c2v_88_out3[QUAN_SIZE-1:0] = c2v_3[88];
assign v2c_3[88] = v2c_88_in3[QUAN_SIZE-1:0];
assign c2v_88_out4[QUAN_SIZE-1:0] = c2v_4[88];
assign v2c_4[88] = v2c_88_in4[QUAN_SIZE-1:0];
assign c2v_88_out5[QUAN_SIZE-1:0] = c2v_5[88];
assign v2c_5[88] = v2c_88_in5[QUAN_SIZE-1:0];
assign c2v_89_out0[QUAN_SIZE-1:0] = c2v_0[89];
assign v2c_0[89] = v2c_89_in0[QUAN_SIZE-1:0];
assign c2v_89_out1[QUAN_SIZE-1:0] = c2v_1[89];
assign v2c_1[89] = v2c_89_in1[QUAN_SIZE-1:0];
assign c2v_89_out2[QUAN_SIZE-1:0] = c2v_2[89];
assign v2c_2[89] = v2c_89_in2[QUAN_SIZE-1:0];
assign c2v_89_out3[QUAN_SIZE-1:0] = c2v_3[89];
assign v2c_3[89] = v2c_89_in3[QUAN_SIZE-1:0];
assign c2v_89_out4[QUAN_SIZE-1:0] = c2v_4[89];
assign v2c_4[89] = v2c_89_in4[QUAN_SIZE-1:0];
assign c2v_89_out5[QUAN_SIZE-1:0] = c2v_5[89];
assign v2c_5[89] = v2c_89_in5[QUAN_SIZE-1:0];
assign c2v_90_out0[QUAN_SIZE-1:0] = c2v_0[90];
assign v2c_0[90] = v2c_90_in0[QUAN_SIZE-1:0];
assign c2v_90_out1[QUAN_SIZE-1:0] = c2v_1[90];
assign v2c_1[90] = v2c_90_in1[QUAN_SIZE-1:0];
assign c2v_90_out2[QUAN_SIZE-1:0] = c2v_2[90];
assign v2c_2[90] = v2c_90_in2[QUAN_SIZE-1:0];
assign c2v_90_out3[QUAN_SIZE-1:0] = c2v_3[90];
assign v2c_3[90] = v2c_90_in3[QUAN_SIZE-1:0];
assign c2v_90_out4[QUAN_SIZE-1:0] = c2v_4[90];
assign v2c_4[90] = v2c_90_in4[QUAN_SIZE-1:0];
assign c2v_90_out5[QUAN_SIZE-1:0] = c2v_5[90];
assign v2c_5[90] = v2c_90_in5[QUAN_SIZE-1:0];
assign c2v_91_out0[QUAN_SIZE-1:0] = c2v_0[91];
assign v2c_0[91] = v2c_91_in0[QUAN_SIZE-1:0];
assign c2v_91_out1[QUAN_SIZE-1:0] = c2v_1[91];
assign v2c_1[91] = v2c_91_in1[QUAN_SIZE-1:0];
assign c2v_91_out2[QUAN_SIZE-1:0] = c2v_2[91];
assign v2c_2[91] = v2c_91_in2[QUAN_SIZE-1:0];
assign c2v_91_out3[QUAN_SIZE-1:0] = c2v_3[91];
assign v2c_3[91] = v2c_91_in3[QUAN_SIZE-1:0];
assign c2v_91_out4[QUAN_SIZE-1:0] = c2v_4[91];
assign v2c_4[91] = v2c_91_in4[QUAN_SIZE-1:0];
assign c2v_91_out5[QUAN_SIZE-1:0] = c2v_5[91];
assign v2c_5[91] = v2c_91_in5[QUAN_SIZE-1:0];
assign c2v_92_out0[QUAN_SIZE-1:0] = c2v_0[92];
assign v2c_0[92] = v2c_92_in0[QUAN_SIZE-1:0];
assign c2v_92_out1[QUAN_SIZE-1:0] = c2v_1[92];
assign v2c_1[92] = v2c_92_in1[QUAN_SIZE-1:0];
assign c2v_92_out2[QUAN_SIZE-1:0] = c2v_2[92];
assign v2c_2[92] = v2c_92_in2[QUAN_SIZE-1:0];
assign c2v_92_out3[QUAN_SIZE-1:0] = c2v_3[92];
assign v2c_3[92] = v2c_92_in3[QUAN_SIZE-1:0];
assign c2v_92_out4[QUAN_SIZE-1:0] = c2v_4[92];
assign v2c_4[92] = v2c_92_in4[QUAN_SIZE-1:0];
assign c2v_92_out5[QUAN_SIZE-1:0] = c2v_5[92];
assign v2c_5[92] = v2c_92_in5[QUAN_SIZE-1:0];
assign c2v_93_out0[QUAN_SIZE-1:0] = c2v_0[93];
assign v2c_0[93] = v2c_93_in0[QUAN_SIZE-1:0];
assign c2v_93_out1[QUAN_SIZE-1:0] = c2v_1[93];
assign v2c_1[93] = v2c_93_in1[QUAN_SIZE-1:0];
assign c2v_93_out2[QUAN_SIZE-1:0] = c2v_2[93];
assign v2c_2[93] = v2c_93_in2[QUAN_SIZE-1:0];
assign c2v_93_out3[QUAN_SIZE-1:0] = c2v_3[93];
assign v2c_3[93] = v2c_93_in3[QUAN_SIZE-1:0];
assign c2v_93_out4[QUAN_SIZE-1:0] = c2v_4[93];
assign v2c_4[93] = v2c_93_in4[QUAN_SIZE-1:0];
assign c2v_93_out5[QUAN_SIZE-1:0] = c2v_5[93];
assign v2c_5[93] = v2c_93_in5[QUAN_SIZE-1:0];
assign c2v_94_out0[QUAN_SIZE-1:0] = c2v_0[94];
assign v2c_0[94] = v2c_94_in0[QUAN_SIZE-1:0];
assign c2v_94_out1[QUAN_SIZE-1:0] = c2v_1[94];
assign v2c_1[94] = v2c_94_in1[QUAN_SIZE-1:0];
assign c2v_94_out2[QUAN_SIZE-1:0] = c2v_2[94];
assign v2c_2[94] = v2c_94_in2[QUAN_SIZE-1:0];
assign c2v_94_out3[QUAN_SIZE-1:0] = c2v_3[94];
assign v2c_3[94] = v2c_94_in3[QUAN_SIZE-1:0];
assign c2v_94_out4[QUAN_SIZE-1:0] = c2v_4[94];
assign v2c_4[94] = v2c_94_in4[QUAN_SIZE-1:0];
assign c2v_94_out5[QUAN_SIZE-1:0] = c2v_5[94];
assign v2c_5[94] = v2c_94_in5[QUAN_SIZE-1:0];
assign c2v_95_out0[QUAN_SIZE-1:0] = c2v_0[95];
assign v2c_0[95] = v2c_95_in0[QUAN_SIZE-1:0];
assign c2v_95_out1[QUAN_SIZE-1:0] = c2v_1[95];
assign v2c_1[95] = v2c_95_in1[QUAN_SIZE-1:0];
assign c2v_95_out2[QUAN_SIZE-1:0] = c2v_2[95];
assign v2c_2[95] = v2c_95_in2[QUAN_SIZE-1:0];
assign c2v_95_out3[QUAN_SIZE-1:0] = c2v_3[95];
assign v2c_3[95] = v2c_95_in3[QUAN_SIZE-1:0];
assign c2v_95_out4[QUAN_SIZE-1:0] = c2v_4[95];
assign v2c_4[95] = v2c_95_in4[QUAN_SIZE-1:0];
assign c2v_95_out5[QUAN_SIZE-1:0] = c2v_5[95];
assign v2c_5[95] = v2c_95_in5[QUAN_SIZE-1:0];
assign c2v_96_out0[QUAN_SIZE-1:0] = c2v_0[96];
assign v2c_0[96] = v2c_96_in0[QUAN_SIZE-1:0];
assign c2v_96_out1[QUAN_SIZE-1:0] = c2v_1[96];
assign v2c_1[96] = v2c_96_in1[QUAN_SIZE-1:0];
assign c2v_96_out2[QUAN_SIZE-1:0] = c2v_2[96];
assign v2c_2[96] = v2c_96_in2[QUAN_SIZE-1:0];
assign c2v_96_out3[QUAN_SIZE-1:0] = c2v_3[96];
assign v2c_3[96] = v2c_96_in3[QUAN_SIZE-1:0];
assign c2v_96_out4[QUAN_SIZE-1:0] = c2v_4[96];
assign v2c_4[96] = v2c_96_in4[QUAN_SIZE-1:0];
assign c2v_96_out5[QUAN_SIZE-1:0] = c2v_5[96];
assign v2c_5[96] = v2c_96_in5[QUAN_SIZE-1:0];
assign c2v_97_out0[QUAN_SIZE-1:0] = c2v_0[97];
assign v2c_0[97] = v2c_97_in0[QUAN_SIZE-1:0];
assign c2v_97_out1[QUAN_SIZE-1:0] = c2v_1[97];
assign v2c_1[97] = v2c_97_in1[QUAN_SIZE-1:0];
assign c2v_97_out2[QUAN_SIZE-1:0] = c2v_2[97];
assign v2c_2[97] = v2c_97_in2[QUAN_SIZE-1:0];
assign c2v_97_out3[QUAN_SIZE-1:0] = c2v_3[97];
assign v2c_3[97] = v2c_97_in3[QUAN_SIZE-1:0];
assign c2v_97_out4[QUAN_SIZE-1:0] = c2v_4[97];
assign v2c_4[97] = v2c_97_in4[QUAN_SIZE-1:0];
assign c2v_97_out5[QUAN_SIZE-1:0] = c2v_5[97];
assign v2c_5[97] = v2c_97_in5[QUAN_SIZE-1:0];
assign c2v_98_out0[QUAN_SIZE-1:0] = c2v_0[98];
assign v2c_0[98] = v2c_98_in0[QUAN_SIZE-1:0];
assign c2v_98_out1[QUAN_SIZE-1:0] = c2v_1[98];
assign v2c_1[98] = v2c_98_in1[QUAN_SIZE-1:0];
assign c2v_98_out2[QUAN_SIZE-1:0] = c2v_2[98];
assign v2c_2[98] = v2c_98_in2[QUAN_SIZE-1:0];
assign c2v_98_out3[QUAN_SIZE-1:0] = c2v_3[98];
assign v2c_3[98] = v2c_98_in3[QUAN_SIZE-1:0];
assign c2v_98_out4[QUAN_SIZE-1:0] = c2v_4[98];
assign v2c_4[98] = v2c_98_in4[QUAN_SIZE-1:0];
assign c2v_98_out5[QUAN_SIZE-1:0] = c2v_5[98];
assign v2c_5[98] = v2c_98_in5[QUAN_SIZE-1:0];
assign c2v_99_out0[QUAN_SIZE-1:0] = c2v_0[99];
assign v2c_0[99] = v2c_99_in0[QUAN_SIZE-1:0];
assign c2v_99_out1[QUAN_SIZE-1:0] = c2v_1[99];
assign v2c_1[99] = v2c_99_in1[QUAN_SIZE-1:0];
assign c2v_99_out2[QUAN_SIZE-1:0] = c2v_2[99];
assign v2c_2[99] = v2c_99_in2[QUAN_SIZE-1:0];
assign c2v_99_out3[QUAN_SIZE-1:0] = c2v_3[99];
assign v2c_3[99] = v2c_99_in3[QUAN_SIZE-1:0];
assign c2v_99_out4[QUAN_SIZE-1:0] = c2v_4[99];
assign v2c_4[99] = v2c_99_in4[QUAN_SIZE-1:0];
assign c2v_99_out5[QUAN_SIZE-1:0] = c2v_5[99];
assign v2c_5[99] = v2c_99_in5[QUAN_SIZE-1:0];
assign c2v_100_out0[QUAN_SIZE-1:0] = c2v_0[100];
assign v2c_0[100] = v2c_100_in0[QUAN_SIZE-1:0];
assign c2v_100_out1[QUAN_SIZE-1:0] = c2v_1[100];
assign v2c_1[100] = v2c_100_in1[QUAN_SIZE-1:0];
assign c2v_100_out2[QUAN_SIZE-1:0] = c2v_2[100];
assign v2c_2[100] = v2c_100_in2[QUAN_SIZE-1:0];
assign c2v_100_out3[QUAN_SIZE-1:0] = c2v_3[100];
assign v2c_3[100] = v2c_100_in3[QUAN_SIZE-1:0];
assign c2v_100_out4[QUAN_SIZE-1:0] = c2v_4[100];
assign v2c_4[100] = v2c_100_in4[QUAN_SIZE-1:0];
assign c2v_100_out5[QUAN_SIZE-1:0] = c2v_5[100];
assign v2c_5[100] = v2c_100_in5[QUAN_SIZE-1:0];
assign c2v_101_out0[QUAN_SIZE-1:0] = c2v_0[101];
assign v2c_0[101] = v2c_101_in0[QUAN_SIZE-1:0];
assign c2v_101_out1[QUAN_SIZE-1:0] = c2v_1[101];
assign v2c_1[101] = v2c_101_in1[QUAN_SIZE-1:0];
assign c2v_101_out2[QUAN_SIZE-1:0] = c2v_2[101];
assign v2c_2[101] = v2c_101_in2[QUAN_SIZE-1:0];
assign c2v_101_out3[QUAN_SIZE-1:0] = c2v_3[101];
assign v2c_3[101] = v2c_101_in3[QUAN_SIZE-1:0];
assign c2v_101_out4[QUAN_SIZE-1:0] = c2v_4[101];
assign v2c_4[101] = v2c_101_in4[QUAN_SIZE-1:0];
assign c2v_101_out5[QUAN_SIZE-1:0] = c2v_5[101];
assign v2c_5[101] = v2c_101_in5[QUAN_SIZE-1:0];
endmodule