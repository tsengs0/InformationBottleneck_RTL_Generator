`define AXI_FRAME_SIZE 32 // the size of one AXI package is 32-bit
`define FRAME_COUNT_SIZE 22