module mem_subsystem_top #(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 85,
	parameter LAYER_NUM = 3,
	// Parameters of extrinsic RAMs
	parameter RAM_UNIT_MSG_NUM = 17, // each RAM unit contributes 17 messages of size 4-bit
	parameter RAM_PORTA_RANGE = 9, // 9 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port A,
	parameter RAM_PORTB_RANGE = 8, // 8 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port b, 
	parameter MEM_DEVICE_NUM = 5,
	parameter DEPTH = 1024,
	parameter WIDTH = 36,
	parameter ADDR = $clog2(DEPTH)
) (
	// The memory Dout port to permutation network for instrinsic messages of variable nodes of upcoming operation
	output wire [QUAN_SIZE-1:0] mem_to_bs_0,
	output wire [QUAN_SIZE-1:0] mem_to_bs_1,
	output wire [QUAN_SIZE-1:0] mem_to_bs_2,
	output wire [QUAN_SIZE-1:0] mem_to_bs_3,
	output wire [QUAN_SIZE-1:0] mem_to_bs_4,
	output wire [QUAN_SIZE-1:0] mem_to_bs_5,
	output wire [QUAN_SIZE-1:0] mem_to_bs_6,
	output wire [QUAN_SIZE-1:0] mem_to_bs_7,
	output wire [QUAN_SIZE-1:0] mem_to_bs_8,
	output wire [QUAN_SIZE-1:0] mem_to_bs_9,
	output wire [QUAN_SIZE-1:0] mem_to_bs_10,
	output wire [QUAN_SIZE-1:0] mem_to_bs_11,
	output wire [QUAN_SIZE-1:0] mem_to_bs_12,
	output wire [QUAN_SIZE-1:0] mem_to_bs_13,
	output wire [QUAN_SIZE-1:0] mem_to_bs_14,
	output wire [QUAN_SIZE-1:0] mem_to_bs_15,
	output wire [QUAN_SIZE-1:0] mem_to_bs_16,
	output wire [QUAN_SIZE-1:0] mem_to_bs_17,
	output wire [QUAN_SIZE-1:0] mem_to_bs_18,
	output wire [QUAN_SIZE-1:0] mem_to_bs_19,
	output wire [QUAN_SIZE-1:0] mem_to_bs_20,
	output wire [QUAN_SIZE-1:0] mem_to_bs_21,
	output wire [QUAN_SIZE-1:0] mem_to_bs_22,
	output wire [QUAN_SIZE-1:0] mem_to_bs_23,
	output wire [QUAN_SIZE-1:0] mem_to_bs_24,
	output wire [QUAN_SIZE-1:0] mem_to_bs_25,
	output wire [QUAN_SIZE-1:0] mem_to_bs_26,
	output wire [QUAN_SIZE-1:0] mem_to_bs_27,
	output wire [QUAN_SIZE-1:0] mem_to_bs_28,
	output wire [QUAN_SIZE-1:0] mem_to_bs_29,
	output wire [QUAN_SIZE-1:0] mem_to_bs_30,
	output wire [QUAN_SIZE-1:0] mem_to_bs_31,
	output wire [QUAN_SIZE-1:0] mem_to_bs_32,
	output wire [QUAN_SIZE-1:0] mem_to_bs_33,
	output wire [QUAN_SIZE-1:0] mem_to_bs_34,
	output wire [QUAN_SIZE-1:0] mem_to_bs_35,
	output wire [QUAN_SIZE-1:0] mem_to_bs_36,
	output wire [QUAN_SIZE-1:0] mem_to_bs_37,
	output wire [QUAN_SIZE-1:0] mem_to_bs_38,
	output wire [QUAN_SIZE-1:0] mem_to_bs_39,
	output wire [QUAN_SIZE-1:0] mem_to_bs_40,
	output wire [QUAN_SIZE-1:0] mem_to_bs_41,
	output wire [QUAN_SIZE-1:0] mem_to_bs_42,
	output wire [QUAN_SIZE-1:0] mem_to_bs_43,
	output wire [QUAN_SIZE-1:0] mem_to_bs_44,
	output wire [QUAN_SIZE-1:0] mem_to_bs_45,
	output wire [QUAN_SIZE-1:0] mem_to_bs_46,
	output wire [QUAN_SIZE-1:0] mem_to_bs_47,
	output wire [QUAN_SIZE-1:0] mem_to_bs_48,
	output wire [QUAN_SIZE-1:0] mem_to_bs_49,
	output wire [QUAN_SIZE-1:0] mem_to_bs_50,
	output wire [QUAN_SIZE-1:0] mem_to_bs_51,
	output wire [QUAN_SIZE-1:0] mem_to_bs_52,
	output wire [QUAN_SIZE-1:0] mem_to_bs_53,
	output wire [QUAN_SIZE-1:0] mem_to_bs_54,
	output wire [QUAN_SIZE-1:0] mem_to_bs_55,
	output wire [QUAN_SIZE-1:0] mem_to_bs_56,
	output wire [QUAN_SIZE-1:0] mem_to_bs_57,
	output wire [QUAN_SIZE-1:0] mem_to_bs_58,
	output wire [QUAN_SIZE-1:0] mem_to_bs_59,
	output wire [QUAN_SIZE-1:0] mem_to_bs_60,
	output wire [QUAN_SIZE-1:0] mem_to_bs_61,
	output wire [QUAN_SIZE-1:0] mem_to_bs_62,
	output wire [QUAN_SIZE-1:0] mem_to_bs_63,
	output wire [QUAN_SIZE-1:0] mem_to_bs_64,
	output wire [QUAN_SIZE-1:0] mem_to_bs_65,
	output wire [QUAN_SIZE-1:0] mem_to_bs_66,
	output wire [QUAN_SIZE-1:0] mem_to_bs_67,
	output wire [QUAN_SIZE-1:0] mem_to_bs_68,
	output wire [QUAN_SIZE-1:0] mem_to_bs_69,
	output wire [QUAN_SIZE-1:0] mem_to_bs_70,
	output wire [QUAN_SIZE-1:0] mem_to_bs_71,
	output wire [QUAN_SIZE-1:0] mem_to_bs_72,
	output wire [QUAN_SIZE-1:0] mem_to_bs_73,
	output wire [QUAN_SIZE-1:0] mem_to_bs_74,
	output wire [QUAN_SIZE-1:0] mem_to_bs_75,
	output wire [QUAN_SIZE-1:0] mem_to_bs_76,
	output wire [QUAN_SIZE-1:0] mem_to_bs_77,
	output wire [QUAN_SIZE-1:0] mem_to_bs_78,
	output wire [QUAN_SIZE-1:0] mem_to_bs_79,
	output wire [QUAN_SIZE-1:0] mem_to_bs_80,
	output wire [QUAN_SIZE-1:0] mem_to_bs_81,
	output wire [QUAN_SIZE-1:0] mem_to_bs_82,
	output wire [QUAN_SIZE-1:0] mem_to_bs_83,
	output wire [QUAN_SIZE-1:0] mem_to_bs_84,
	// The memory Dout port to check nodes as instrinsic messages
	output wire [QUAN_SIZE-1:0] mem_to_cnu_0,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_1,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_2,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_3,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_4,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_5,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_6,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_7,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_8,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_9,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_10,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_11,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_12,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_13,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_14,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_15,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_16,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_17,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_18,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_19,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_20,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_21,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_22,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_23,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_24,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_25,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_26,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_27,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_28,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_29,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_30,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_31,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_32,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_33,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_34,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_35,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_36,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_37,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_38,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_39,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_40,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_41,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_42,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_43,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_44,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_45,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_46,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_47,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_48,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_49,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_50,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_51,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_52,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_53,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_54,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_55,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_56,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_57,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_58,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_59,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_60,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_61,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_62,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_63,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_64,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_65,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_66,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_67,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_68,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_69,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_70,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_71,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_72,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_73,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_74,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_75,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_76,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_77,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_78,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_79,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_80,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_81,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_82,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_83,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_84,

	input wire [QUAN_SIZE-1:0] vnu_to_mem_1,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_1,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_2,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_3,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_4,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_5,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_6,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_7,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_8,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_9,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_10,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_11,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_12,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_13,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_14,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_15,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_16,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_17,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_18,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_19,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_20,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_21,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_22,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_23,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_24,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_25,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_26,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_27,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_28,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_29,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_30,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_31,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_32,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_33,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_34,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_35,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_36,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_37,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_38,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_39,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_40,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_41,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_42,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_43,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_44,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_45,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_46,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_47,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_48,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_49,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_50,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_51,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_52,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_53,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_54,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_55,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_56,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_57,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_58,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_59,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_60,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_61,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_62,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_63,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_64,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_65,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_66,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_67,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_68,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_69,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_70,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_71,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_72,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_73,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_74,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_75,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_76,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_77,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_78,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_79,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_80,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_81,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_82,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_83,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_84,

	input wire [QUAN_SIZE-1:0] cnu_to_mem_0,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_1,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_2,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_3,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_4,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_5,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_6,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_7,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_8,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_9,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_10,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_11,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_12,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_13,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_14,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_15,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_16,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_17,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_18,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_19,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_20,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_21,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_22,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_23,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_24,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_25,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_26,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_27,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_28,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_29,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_30,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_31,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_32,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_33,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_34,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_35,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_36,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_37,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_38,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_39,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_40,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_41,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_42,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_43,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_44,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_45,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_46,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_47,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_48,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_49,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_50,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_51,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_52,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_53,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_54,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_55,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_56,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_57,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_58,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_59,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_60,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_61,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_62,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_63,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_64,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_65,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_66,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_67,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_68,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_69,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_70,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_71,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_72,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_73,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_74,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_75,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_76,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_77,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_78,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_79,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_80,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_81,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_82,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_83,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_84,

	input wire sched_cmd, // 1'b0: align_in from variable msg; 1'b1: align_in from check msg
	input wire [CHECK_PARALLELISM-1:0] delay_cmd,
	input wire [ADDR-1:0] sync_addr,
	input wire [LAYER_NUM-1:0] layer_status,
	input wire first_row_chunk,
	input wire we,
	input wire sys_clk,
	input wire rstn
);

// Memory Input Interface where page-aligned mechanism is embedded insight
wire [QUAN_SIZE-1:0] page_align_out [0:CHECK_PARALLELISM-1];
ram_pageAlign_interface #(
	.QUAN_SIZE (QUAN_SIZE), //4
	.CHECK_PARALLELISM (CHECK_PARALLELISM), // 85
	.LAYER_NUM (LAYER_NUM) // 3
) ram_pageAlign_interface_u0 (
	.msg_out_0  (page_align_out[0 ]),
	.msg_out_1  (page_align_out[1 ]),
	.msg_out_2  (page_align_out[2 ]),
	.msg_out_3  (page_align_out[3 ]),
	.msg_out_4  (page_align_out[4 ]),
	.msg_out_5  (page_align_out[5 ]),
	.msg_out_6  (page_align_out[6 ]),
	.msg_out_7  (page_align_out[7 ]),
	.msg_out_8  (page_align_out[8 ]),
	.msg_out_9  (page_align_out[9 ]),
	.msg_out_10 (page_align_out[10]),
	.msg_out_11 (page_align_out[11]),
	.msg_out_12 (page_align_out[12]),
	.msg_out_13 (page_align_out[13]),
	.msg_out_14 (page_align_out[14]),
	.msg_out_15 (page_align_out[15]),
	.msg_out_16 (page_align_out[16]),
	.msg_out_17 (page_align_out[17]),
	.msg_out_18 (page_align_out[18]),
	.msg_out_19 (page_align_out[19]),
	.msg_out_20 (page_align_out[20]),
	.msg_out_21 (page_align_out[21]),
	.msg_out_22 (page_align_out[22]),
	.msg_out_23 (page_align_out[23]),
	.msg_out_24 (page_align_out[24]),
	.msg_out_25 (page_align_out[25]),
	.msg_out_26 (page_align_out[26]),
	.msg_out_27 (page_align_out[27]),
	.msg_out_28 (page_align_out[28]),
	.msg_out_29 (page_align_out[29]),
	.msg_out_30 (page_align_out[30]),
	.msg_out_31 (page_align_out[31]),
	.msg_out_32 (page_align_out[32]),
	.msg_out_33 (page_align_out[33]),
	.msg_out_34 (page_align_out[34]),
	.msg_out_35 (page_align_out[35]),
	.msg_out_36 (page_align_out[36]),
	.msg_out_37 (page_align_out[37]),
	.msg_out_38 (page_align_out[38]),
	.msg_out_39 (page_align_out[39]),
	.msg_out_40 (page_align_out[40]),
	.msg_out_41 (page_align_out[41]),
	.msg_out_42 (page_align_out[42]),
	.msg_out_43 (page_align_out[43]),
	.msg_out_44 (page_align_out[44]),
	.msg_out_45 (page_align_out[45]),
	.msg_out_46 (page_align_out[46]),
	.msg_out_47 (page_align_out[47]),
	.msg_out_48 (page_align_out[48]),
	.msg_out_49 (page_align_out[49]),
	.msg_out_50 (page_align_out[50]),
	.msg_out_51 (page_align_out[51]),
	.msg_out_52 (page_align_out[52]),
	.msg_out_53 (page_align_out[53]),
	.msg_out_54 (page_align_out[54]),
	.msg_out_55 (page_align_out[55]),
	.msg_out_56 (page_align_out[56]),
	.msg_out_57 (page_align_out[57]),
	.msg_out_58 (page_align_out[58]),
	.msg_out_59 (page_align_out[59]),
	.msg_out_60 (page_align_out[60]),
	.msg_out_61 (page_align_out[61]),
	.msg_out_62 (page_align_out[62]),
	.msg_out_63 (page_align_out[63]),
	.msg_out_64 (page_align_out[64]),
	.msg_out_65 (page_align_out[65]),
	.msg_out_66 (page_align_out[66]),
	.msg_out_67 (page_align_out[67]),
	.msg_out_68 (page_align_out[68]),
	.msg_out_69 (page_align_out[69]),
	.msg_out_70 (page_align_out[70]),
	.msg_out_71 (page_align_out[71]),
	.msg_out_72 (page_align_out[72]),
	.msg_out_73 (page_align_out[73]),
	.msg_out_74 (page_align_out[74]),
	.msg_out_75 (page_align_out[75]),
	.msg_out_76 (page_align_out[76]),
	.msg_out_77 (page_align_out[77]),
	.msg_out_78 (page_align_out[78]),
	.msg_out_79 (page_align_out[79]),
	.msg_out_80 (page_align_out[80]),
	.msg_out_81 (page_align_out[81]),
	.msg_out_82 (page_align_out[82]),
	.msg_out_83 (page_align_out[83]),
	.msg_out_84 (page_align_out[84]),

	.vnu_msg_in_0  (vnu_to_mem_1 [QUAN_SIZE-1:0]),
	.vnu_msg_in_1  (vnu_to_mem_1 [QUAN_SIZE-1:0]),
	.vnu_msg_in_2  (vnu_to_mem_2 [QUAN_SIZE-1:0]),
	.vnu_msg_in_3  (vnu_to_mem_3 [QUAN_SIZE-1:0]),
	.vnu_msg_in_4  (vnu_to_mem_4 [QUAN_SIZE-1:0]),
	.vnu_msg_in_5  (vnu_to_mem_5 [QUAN_SIZE-1:0]),
	.vnu_msg_in_6  (vnu_to_mem_6 [QUAN_SIZE-1:0]),
	.vnu_msg_in_7  (vnu_to_mem_7 [QUAN_SIZE-1:0]),
	.vnu_msg_in_8  (vnu_to_mem_8 [QUAN_SIZE-1:0]),
	.vnu_msg_in_9  (vnu_to_mem_9 [QUAN_SIZE-1:0]),
	.vnu_msg_in_10 (vnu_to_mem_10[QUAN_SIZE-1:0]),
	.vnu_msg_in_11 (vnu_to_mem_11[QUAN_SIZE-1:0]),
	.vnu_msg_in_12 (vnu_to_mem_12[QUAN_SIZE-1:0]),
	.vnu_msg_in_13 (vnu_to_mem_13[QUAN_SIZE-1:0]),
	.vnu_msg_in_14 (vnu_to_mem_14[QUAN_SIZE-1:0]),
	.vnu_msg_in_15 (vnu_to_mem_15[QUAN_SIZE-1:0]),
	.vnu_msg_in_16 (vnu_to_mem_16[QUAN_SIZE-1:0]),
	.vnu_msg_in_17 (vnu_to_mem_17[QUAN_SIZE-1:0]),
	.vnu_msg_in_18 (vnu_to_mem_18[QUAN_SIZE-1:0]),
	.vnu_msg_in_19 (vnu_to_mem_19[QUAN_SIZE-1:0]),
	.vnu_msg_in_20 (vnu_to_mem_20[QUAN_SIZE-1:0]),
	.vnu_msg_in_21 (vnu_to_mem_21[QUAN_SIZE-1:0]),
	.vnu_msg_in_22 (vnu_to_mem_22[QUAN_SIZE-1:0]),
	.vnu_msg_in_23 (vnu_to_mem_23[QUAN_SIZE-1:0]),
	.vnu_msg_in_24 (vnu_to_mem_24[QUAN_SIZE-1:0]),
	.vnu_msg_in_25 (vnu_to_mem_25[QUAN_SIZE-1:0]),
	.vnu_msg_in_26 (vnu_to_mem_26[QUAN_SIZE-1:0]),
	.vnu_msg_in_27 (vnu_to_mem_27[QUAN_SIZE-1:0]),
	.vnu_msg_in_28 (vnu_to_mem_28[QUAN_SIZE-1:0]),
	.vnu_msg_in_29 (vnu_to_mem_29[QUAN_SIZE-1:0]),
	.vnu_msg_in_30 (vnu_to_mem_30[QUAN_SIZE-1:0]),
	.vnu_msg_in_31 (vnu_to_mem_31[QUAN_SIZE-1:0]),
	.vnu_msg_in_32 (vnu_to_mem_32[QUAN_SIZE-1:0]),
	.vnu_msg_in_33 (vnu_to_mem_33[QUAN_SIZE-1:0]),
	.vnu_msg_in_34 (vnu_to_mem_34[QUAN_SIZE-1:0]),
	.vnu_msg_in_35 (vnu_to_mem_35[QUAN_SIZE-1:0]),
	.vnu_msg_in_36 (vnu_to_mem_36[QUAN_SIZE-1:0]),
	.vnu_msg_in_37 (vnu_to_mem_37[QUAN_SIZE-1:0]),
	.vnu_msg_in_38 (vnu_to_mem_38[QUAN_SIZE-1:0]),
	.vnu_msg_in_39 (vnu_to_mem_39[QUAN_SIZE-1:0]),
	.vnu_msg_in_40 (vnu_to_mem_40[QUAN_SIZE-1:0]),
	.vnu_msg_in_41 (vnu_to_mem_41[QUAN_SIZE-1:0]),
	.vnu_msg_in_42 (vnu_to_mem_42[QUAN_SIZE-1:0]),
	.vnu_msg_in_43 (vnu_to_mem_43[QUAN_SIZE-1:0]),
	.vnu_msg_in_44 (vnu_to_mem_44[QUAN_SIZE-1:0]),
	.vnu_msg_in_45 (vnu_to_mem_45[QUAN_SIZE-1:0]),
	.vnu_msg_in_46 (vnu_to_mem_46[QUAN_SIZE-1:0]),
	.vnu_msg_in_47 (vnu_to_mem_47[QUAN_SIZE-1:0]),
	.vnu_msg_in_48 (vnu_to_mem_48[QUAN_SIZE-1:0]),
	.vnu_msg_in_49 (vnu_to_mem_49[QUAN_SIZE-1:0]),
	.vnu_msg_in_50 (vnu_to_mem_50[QUAN_SIZE-1:0]),
	.vnu_msg_in_51 (vnu_to_mem_51[QUAN_SIZE-1:0]),
	.vnu_msg_in_52 (vnu_to_mem_52[QUAN_SIZE-1:0]),
	.vnu_msg_in_53 (vnu_to_mem_53[QUAN_SIZE-1:0]),
	.vnu_msg_in_54 (vnu_to_mem_54[QUAN_SIZE-1:0]),
	.vnu_msg_in_55 (vnu_to_mem_55[QUAN_SIZE-1:0]),
	.vnu_msg_in_56 (vnu_to_mem_56[QUAN_SIZE-1:0]),
	.vnu_msg_in_57 (vnu_to_mem_57[QUAN_SIZE-1:0]),
	.vnu_msg_in_58 (vnu_to_mem_58[QUAN_SIZE-1:0]),
	.vnu_msg_in_59 (vnu_to_mem_59[QUAN_SIZE-1:0]),
	.vnu_msg_in_60 (vnu_to_mem_60[QUAN_SIZE-1:0]),
	.vnu_msg_in_61 (vnu_to_mem_61[QUAN_SIZE-1:0]),
	.vnu_msg_in_62 (vnu_to_mem_62[QUAN_SIZE-1:0]),
	.vnu_msg_in_63 (vnu_to_mem_63[QUAN_SIZE-1:0]),
	.vnu_msg_in_64 (vnu_to_mem_64[QUAN_SIZE-1:0]),
	.vnu_msg_in_65 (vnu_to_mem_65[QUAN_SIZE-1:0]),
	.vnu_msg_in_66 (vnu_to_mem_66[QUAN_SIZE-1:0]),
	.vnu_msg_in_67 (vnu_to_mem_67[QUAN_SIZE-1:0]),
	.vnu_msg_in_68 (vnu_to_mem_68[QUAN_SIZE-1:0]),
	.vnu_msg_in_69 (vnu_to_mem_69[QUAN_SIZE-1:0]),
	.vnu_msg_in_70 (vnu_to_mem_70[QUAN_SIZE-1:0]),
	.vnu_msg_in_71 (vnu_to_mem_71[QUAN_SIZE-1:0]),
	.vnu_msg_in_72 (vnu_to_mem_72[QUAN_SIZE-1:0]),
	.vnu_msg_in_73 (vnu_to_mem_73[QUAN_SIZE-1:0]),
	.vnu_msg_in_74 (vnu_to_mem_74[QUAN_SIZE-1:0]),
	.vnu_msg_in_75 (vnu_to_mem_75[QUAN_SIZE-1:0]),
	.vnu_msg_in_76 (vnu_to_mem_76[QUAN_SIZE-1:0]),
	.vnu_msg_in_77 (vnu_to_mem_77[QUAN_SIZE-1:0]),
	.vnu_msg_in_78 (vnu_to_mem_78[QUAN_SIZE-1:0]),
	.vnu_msg_in_79 (vnu_to_mem_79[QUAN_SIZE-1:0]),
	.vnu_msg_in_80 (vnu_to_mem_80[QUAN_SIZE-1:0]),
	.vnu_msg_in_81 (vnu_to_mem_81[QUAN_SIZE-1:0]),
	.vnu_msg_in_82 (vnu_to_mem_82[QUAN_SIZE-1:0]),
	.vnu_msg_in_83 (vnu_to_mem_83[QUAN_SIZE-1:0]),
	.vnu_msg_in_84 (vnu_to_mem_84[QUAN_SIZE-1:0]),

	.cnu_msg_in_0  (cnu_to_mem_0 [QUAN_SIZE-1:0]),
	.cnu_msg_in_1  (cnu_to_mem_1 [QUAN_SIZE-1:0]),
	.cnu_msg_in_2  (cnu_to_mem_2 [QUAN_SIZE-1:0]),
	.cnu_msg_in_3  (cnu_to_mem_3 [QUAN_SIZE-1:0]),
	.cnu_msg_in_4  (cnu_to_mem_4 [QUAN_SIZE-1:0]),
	.cnu_msg_in_5  (cnu_to_mem_5 [QUAN_SIZE-1:0]),
	.cnu_msg_in_6  (cnu_to_mem_6 [QUAN_SIZE-1:0]),
	.cnu_msg_in_7  (cnu_to_mem_7 [QUAN_SIZE-1:0]),
	.cnu_msg_in_8  (cnu_to_mem_8 [QUAN_SIZE-1:0]),
	.cnu_msg_in_9  (cnu_to_mem_9 [QUAN_SIZE-1:0]),
	.cnu_msg_in_10 (cnu_to_mem_10[QUAN_SIZE-1:0]),
	.cnu_msg_in_11 (cnu_to_mem_11[QUAN_SIZE-1:0]),
	.cnu_msg_in_12 (cnu_to_mem_12[QUAN_SIZE-1:0]),
	.cnu_msg_in_13 (cnu_to_mem_13[QUAN_SIZE-1:0]),
	.cnu_msg_in_14 (cnu_to_mem_14[QUAN_SIZE-1:0]),
	.cnu_msg_in_15 (cnu_to_mem_15[QUAN_SIZE-1:0]),
	.cnu_msg_in_16 (cnu_to_mem_16[QUAN_SIZE-1:0]),
	.cnu_msg_in_17 (cnu_to_mem_17[QUAN_SIZE-1:0]),
	.cnu_msg_in_18 (cnu_to_mem_18[QUAN_SIZE-1:0]),
	.cnu_msg_in_19 (cnu_to_mem_19[QUAN_SIZE-1:0]),
	.cnu_msg_in_20 (cnu_to_mem_20[QUAN_SIZE-1:0]),
	.cnu_msg_in_21 (cnu_to_mem_21[QUAN_SIZE-1:0]),
	.cnu_msg_in_22 (cnu_to_mem_22[QUAN_SIZE-1:0]),
	.cnu_msg_in_23 (cnu_to_mem_23[QUAN_SIZE-1:0]),
	.cnu_msg_in_24 (cnu_to_mem_24[QUAN_SIZE-1:0]),
	.cnu_msg_in_25 (cnu_to_mem_25[QUAN_SIZE-1:0]),
	.cnu_msg_in_26 (cnu_to_mem_26[QUAN_SIZE-1:0]),
	.cnu_msg_in_27 (cnu_to_mem_27[QUAN_SIZE-1:0]),
	.cnu_msg_in_28 (cnu_to_mem_28[QUAN_SIZE-1:0]),
	.cnu_msg_in_29 (cnu_to_mem_29[QUAN_SIZE-1:0]),
	.cnu_msg_in_30 (cnu_to_mem_30[QUAN_SIZE-1:0]),
	.cnu_msg_in_31 (cnu_to_mem_31[QUAN_SIZE-1:0]),
	.cnu_msg_in_32 (cnu_to_mem_32[QUAN_SIZE-1:0]),
	.cnu_msg_in_33 (cnu_to_mem_33[QUAN_SIZE-1:0]),
	.cnu_msg_in_34 (cnu_to_mem_34[QUAN_SIZE-1:0]),
	.cnu_msg_in_35 (cnu_to_mem_35[QUAN_SIZE-1:0]),
	.cnu_msg_in_36 (cnu_to_mem_36[QUAN_SIZE-1:0]),
	.cnu_msg_in_37 (cnu_to_mem_37[QUAN_SIZE-1:0]),
	.cnu_msg_in_38 (cnu_to_mem_38[QUAN_SIZE-1:0]),
	.cnu_msg_in_39 (cnu_to_mem_39[QUAN_SIZE-1:0]),
	.cnu_msg_in_40 (cnu_to_mem_40[QUAN_SIZE-1:0]),
	.cnu_msg_in_41 (cnu_to_mem_41[QUAN_SIZE-1:0]),
	.cnu_msg_in_42 (cnu_to_mem_42[QUAN_SIZE-1:0]),
	.cnu_msg_in_43 (cnu_to_mem_43[QUAN_SIZE-1:0]),
	.cnu_msg_in_44 (cnu_to_mem_44[QUAN_SIZE-1:0]),
	.cnu_msg_in_45 (cnu_to_mem_45[QUAN_SIZE-1:0]),
	.cnu_msg_in_46 (cnu_to_mem_46[QUAN_SIZE-1:0]),
	.cnu_msg_in_47 (cnu_to_mem_47[QUAN_SIZE-1:0]),
	.cnu_msg_in_48 (cnu_to_mem_48[QUAN_SIZE-1:0]),
	.cnu_msg_in_49 (cnu_to_mem_49[QUAN_SIZE-1:0]),
	.cnu_msg_in_50 (cnu_to_mem_50[QUAN_SIZE-1:0]),
	.cnu_msg_in_51 (cnu_to_mem_51[QUAN_SIZE-1:0]),
	.cnu_msg_in_52 (cnu_to_mem_52[QUAN_SIZE-1:0]),
	.cnu_msg_in_53 (cnu_to_mem_53[QUAN_SIZE-1:0]),
	.cnu_msg_in_54 (cnu_to_mem_54[QUAN_SIZE-1:0]),
	.cnu_msg_in_55 (cnu_to_mem_55[QUAN_SIZE-1:0]),
	.cnu_msg_in_56 (cnu_to_mem_56[QUAN_SIZE-1:0]),
	.cnu_msg_in_57 (cnu_to_mem_57[QUAN_SIZE-1:0]),
	.cnu_msg_in_58 (cnu_to_mem_58[QUAN_SIZE-1:0]),
	.cnu_msg_in_59 (cnu_to_mem_59[QUAN_SIZE-1:0]),
	.cnu_msg_in_60 (cnu_to_mem_60[QUAN_SIZE-1:0]),
	.cnu_msg_in_61 (cnu_to_mem_61[QUAN_SIZE-1:0]),
	.cnu_msg_in_62 (cnu_to_mem_62[QUAN_SIZE-1:0]),
	.cnu_msg_in_63 (cnu_to_mem_63[QUAN_SIZE-1:0]),
	.cnu_msg_in_64 (cnu_to_mem_64[QUAN_SIZE-1:0]),
	.cnu_msg_in_65 (cnu_to_mem_65[QUAN_SIZE-1:0]),
	.cnu_msg_in_66 (cnu_to_mem_66[QUAN_SIZE-1:0]),
	.cnu_msg_in_67 (cnu_to_mem_67[QUAN_SIZE-1:0]),
	.cnu_msg_in_68 (cnu_to_mem_68[QUAN_SIZE-1:0]),
	.cnu_msg_in_69 (cnu_to_mem_69[QUAN_SIZE-1:0]),
	.cnu_msg_in_70 (cnu_to_mem_70[QUAN_SIZE-1:0]),
	.cnu_msg_in_71 (cnu_to_mem_71[QUAN_SIZE-1:0]),
	.cnu_msg_in_72 (cnu_to_mem_72[QUAN_SIZE-1:0]),
	.cnu_msg_in_73 (cnu_to_mem_73[QUAN_SIZE-1:0]),
	.cnu_msg_in_74 (cnu_to_mem_74[QUAN_SIZE-1:0]),
	.cnu_msg_in_75 (cnu_to_mem_75[QUAN_SIZE-1:0]),
	.cnu_msg_in_76 (cnu_to_mem_76[QUAN_SIZE-1:0]),
	.cnu_msg_in_77 (cnu_to_mem_77[QUAN_SIZE-1:0]),
	.cnu_msg_in_78 (cnu_to_mem_78[QUAN_SIZE-1:0]),
	.cnu_msg_in_79 (cnu_to_mem_79[QUAN_SIZE-1:0]),
	.cnu_msg_in_80 (cnu_to_mem_80[QUAN_SIZE-1:0]),
	.cnu_msg_in_81 (cnu_to_mem_81[QUAN_SIZE-1:0]),
	.cnu_msg_in_82 (cnu_to_mem_82[QUAN_SIZE-1:0]),
	.cnu_msg_in_83 (cnu_to_mem_83[QUAN_SIZE-1:0]),
	.cnu_msg_in_84 (cnu_to_mem_84[QUAN_SIZE-1:0]),

	.sched_cmd (sched_cmd), // 1'b0: align_in from variable msg; 1'b1: align_in from check msg
	.delay_cmd (delay_cmd[CHECK_PARALLELISM-1:0]),
	.layer_status (layer_status[LAYER_NUM-1:0]),
	.first_row_chunk (first_row_chunk),
	.sys_clk (sys_clk),
	.rstn (rstn)
);

// Extrinsic RAM instatiation
wire [QUAN_SIZE-1:0] ram_dout_reg [0:CHECK_PARALLELISM-1];
column_ram_pc85 #(
	.QUAN_SIZE(QUAN_SIZE),
	.CHECK_PARALLELISM(CHECK_PARALLELISM),
	.RAM_UNIT_MSG_NUM(RAM_UNIT_MSG_NUM),
	.RAM_PORTA_RANGE(RAM_PORTA_RANGE),
	.RAM_PORTB_RANGE(RAM_PORTB_RANGE),
	.MEM_DEVICE_NUM(MEM_DEVICE_NUM),
	.DEPTH(DEPTH),
	.WIDTH(WIDTH),
	.ADDR(ADDR)
) inst_column_ram_pc85 (
	.Dout_0    (ram_dout_reg[0 ]),
	.Dout_1    (ram_dout_reg[1 ]),
	.Dout_2    (ram_dout_reg[2 ]),
	.Dout_3    (ram_dout_reg[3 ]),
	.Dout_4    (ram_dout_reg[4 ]),
	.Dout_5    (ram_dout_reg[5 ]),
	.Dout_6    (ram_dout_reg[6 ]),
	.Dout_7    (ram_dout_reg[7 ]),
	.Dout_8    (ram_dout_reg[8 ]),
	.Dout_9    (ram_dout_reg[9 ]),
	.Dout_10   (ram_dout_reg[10]),
	.Dout_11   (ram_dout_reg[11]),
	.Dout_12   (ram_dout_reg[12]),
	.Dout_13   (ram_dout_reg[13]),
	.Dout_14   (ram_dout_reg[14]),
	.Dout_15   (ram_dout_reg[15]),
	.Dout_16   (ram_dout_reg[16]),
	.Dout_17   (ram_dout_reg[17]),
	.Dout_18   (ram_dout_reg[18]),
	.Dout_19   (ram_dout_reg[19]),
	.Dout_20   (ram_dout_reg[20]),
	.Dout_21   (ram_dout_reg[21]),
	.Dout_22   (ram_dout_reg[22]),
	.Dout_23   (ram_dout_reg[23]),
	.Dout_24   (ram_dout_reg[24]),
	.Dout_25   (ram_dout_reg[25]),
	.Dout_26   (ram_dout_reg[26]),
	.Dout_27   (ram_dout_reg[27]),
	.Dout_28   (ram_dout_reg[28]),
	.Dout_29   (ram_dout_reg[29]),
	.Dout_30   (ram_dout_reg[30]),
	.Dout_31   (ram_dout_reg[31]),
	.Dout_32   (ram_dout_reg[32]),
	.Dout_33   (ram_dout_reg[33]),
	.Dout_34   (ram_dout_reg[34]),
	.Dout_35   (ram_dout_reg[35]),
	.Dout_36   (ram_dout_reg[36]),
	.Dout_37   (ram_dout_reg[37]),
	.Dout_38   (ram_dout_reg[38]),
	.Dout_39   (ram_dout_reg[39]),
	.Dout_40   (ram_dout_reg[40]),
	.Dout_41   (ram_dout_reg[41]),
	.Dout_42   (ram_dout_reg[42]),
	.Dout_43   (ram_dout_reg[43]),
	.Dout_44   (ram_dout_reg[44]),
	.Dout_45   (ram_dout_reg[45]),
	.Dout_46   (ram_dout_reg[46]),
	.Dout_47   (ram_dout_reg[47]),
	.Dout_48   (ram_dout_reg[48]),
	.Dout_49   (ram_dout_reg[49]),
	.Dout_50   (ram_dout_reg[50]),
	.Dout_51   (ram_dout_reg[51]),
	.Dout_52   (ram_dout_reg[52]),
	.Dout_53   (ram_dout_reg[53]),
	.Dout_54   (ram_dout_reg[54]),
	.Dout_55   (ram_dout_reg[55]),
	.Dout_56   (ram_dout_reg[56]),
	.Dout_57   (ram_dout_reg[57]),
	.Dout_58   (ram_dout_reg[58]),
	.Dout_59   (ram_dout_reg[59]),
	.Dout_60   (ram_dout_reg[60]),
	.Dout_61   (ram_dout_reg[61]),
	.Dout_62   (ram_dout_reg[62]),
	.Dout_63   (ram_dout_reg[63]),
	.Dout_64   (ram_dout_reg[64]),
	.Dout_65   (ram_dout_reg[65]),
	.Dout_66   (ram_dout_reg[66]),
	.Dout_67   (ram_dout_reg[67]),
	.Dout_68   (ram_dout_reg[68]),
	.Dout_69   (ram_dout_reg[69]),
	.Dout_70   (ram_dout_reg[70]),
	.Dout_71   (ram_dout_reg[71]),
	.Dout_72   (ram_dout_reg[72]),
	.Dout_73   (ram_dout_reg[73]),
	.Dout_74   (ram_dout_reg[74]),
	.Dout_75   (ram_dout_reg[75]),
	.Dout_76   (ram_dout_reg[76]),
	.Dout_77   (ram_dout_reg[77]),
	.Dout_78   (ram_dout_reg[78]),
	.Dout_79   (ram_dout_reg[79]),
	.Dout_80   (ram_dout_reg[80]),
	.Dout_81   (ram_dout_reg[81]),
	.Dout_82   (ram_dout_reg[82]),
	.Dout_83   (ram_dout_reg[83]),
	.Dout_84   (ram_dout_reg[84]),

	.Din_0     (page_align_out[0 ]),
	.Din_1     (page_align_out[1 ]),
	.Din_2     (page_align_out[2 ]),
	.Din_3     (page_align_out[3 ]),
	.Din_4     (page_align_out[4 ]),
	.Din_5     (page_align_out[5 ]),
	.Din_6     (page_align_out[6 ]),
	.Din_7     (page_align_out[7 ]),
	.Din_8     (page_align_out[8 ]),
	.Din_9     (page_align_out[9 ]),
	.Din_10    (page_align_out[10]),
	.Din_11    (page_align_out[11]),
	.Din_12    (page_align_out[12]),
	.Din_13    (page_align_out[13]),
	.Din_14    (page_align_out[14]),
	.Din_15    (page_align_out[15]),
	.Din_16    (page_align_out[16]),
	.Din_17    (page_align_out[17]),
	.Din_18    (page_align_out[18]),
	.Din_19    (page_align_out[19]),
	.Din_20    (page_align_out[20]),
	.Din_21    (page_align_out[21]),
	.Din_22    (page_align_out[22]),
	.Din_23    (page_align_out[23]),
	.Din_24    (page_align_out[24]),
	.Din_25    (page_align_out[25]),
	.Din_26    (page_align_out[26]),
	.Din_27    (page_align_out[27]),
	.Din_28    (page_align_out[28]),
	.Din_29    (page_align_out[29]),
	.Din_30    (page_align_out[30]),
	.Din_31    (page_align_out[31]),
	.Din_32    (page_align_out[32]),
	.Din_33    (page_align_out[33]),
	.Din_34    (page_align_out[34]),
	.Din_35    (page_align_out[35]),
	.Din_36    (page_align_out[36]),
	.Din_37    (page_align_out[37]),
	.Din_38    (page_align_out[38]),
	.Din_39    (page_align_out[39]),
	.Din_40    (page_align_out[40]),
	.Din_41    (page_align_out[41]),
	.Din_42    (page_align_out[42]),
	.Din_43    (page_align_out[43]),
	.Din_44    (page_align_out[44]),
	.Din_45    (page_align_out[45]),
	.Din_46    (page_align_out[46]),
	.Din_47    (page_align_out[47]),
	.Din_48    (page_align_out[48]),
	.Din_49    (page_align_out[49]),
	.Din_50    (page_align_out[50]),
	.Din_51    (page_align_out[51]),
	.Din_52    (page_align_out[52]),
	.Din_53    (page_align_out[53]),
	.Din_54    (page_align_out[54]),
	.Din_55    (page_align_out[55]),
	.Din_56    (page_align_out[56]),
	.Din_57    (page_align_out[57]),
	.Din_58    (page_align_out[58]),
	.Din_59    (page_align_out[59]),
	.Din_60    (page_align_out[60]),
	.Din_61    (page_align_out[61]),
	.Din_62    (page_align_out[62]),
	.Din_63    (page_align_out[63]),
	.Din_64    (page_align_out[64]),
	.Din_65    (page_align_out[65]),
	.Din_66    (page_align_out[66]),
	.Din_67    (page_align_out[67]),
	.Din_68    (page_align_out[68]),
	.Din_69    (page_align_out[69]),
	.Din_70    (page_align_out[70]),
	.Din_71    (page_align_out[71]),
	.Din_72    (page_align_out[72]),
	.Din_73    (page_align_out[73]),
	.Din_74    (page_align_out[74]),
	.Din_75    (page_align_out[75]),
	.Din_76    (page_align_out[76]),
	.Din_77    (page_align_out[77]),
	.Din_78    (page_align_out[78]),
	.Din_79    (page_align_out[79]),
	.Din_80    (page_align_out[80]),
	.Din_81    (page_align_out[81]),
	.Din_82    (page_align_out[82]),
	.Din_83    (page_align_out[83]),
	.Din_84    (page_align_out[84]),

	.sync_addr (sync_addr),
	.we        (we),
	.sys_clk   (sys_clk)
);

// Final output port - De-multiplexers to either:
// 1) permutation network (outgoing to VNUs) or
// 2) CNUs as instrinsic messages
ram_out_demux #(
	.QUAN_SIZE (QUAN_SIZE), //4
	.CHECK_PARALLELISM (CHECK_PARALLELISM) //85
) ram_out_demux_u0 (
	// The memory Dout port to permutation network for instrinsic messages of variable nodes of upcoming operation
	.mem_to_bs_0  (mem_to_bs_0 ),
	.mem_to_bs_1  (mem_to_bs_1 ),
	.mem_to_bs_2  (mem_to_bs_2 ),
	.mem_to_bs_3  (mem_to_bs_3 ),
	.mem_to_bs_4  (mem_to_bs_4 ),
	.mem_to_bs_5  (mem_to_bs_5 ),
	.mem_to_bs_6  (mem_to_bs_6 ),
	.mem_to_bs_7  (mem_to_bs_7 ),
	.mem_to_bs_8  (mem_to_bs_8 ),
	.mem_to_bs_9  (mem_to_bs_9 ),
	.mem_to_bs_10 (mem_to_bs_10),
	.mem_to_bs_11 (mem_to_bs_11),
	.mem_to_bs_12 (mem_to_bs_12),
	.mem_to_bs_13 (mem_to_bs_13),
	.mem_to_bs_14 (mem_to_bs_14),
	.mem_to_bs_15 (mem_to_bs_15),
	.mem_to_bs_16 (mem_to_bs_16),
	.mem_to_bs_17 (mem_to_bs_17),
	.mem_to_bs_18 (mem_to_bs_18),
	.mem_to_bs_19 (mem_to_bs_19),
	.mem_to_bs_20 (mem_to_bs_20),
	.mem_to_bs_21 (mem_to_bs_21),
	.mem_to_bs_22 (mem_to_bs_22),
	.mem_to_bs_23 (mem_to_bs_23),
	.mem_to_bs_24 (mem_to_bs_24),
	.mem_to_bs_25 (mem_to_bs_25),
	.mem_to_bs_26 (mem_to_bs_26),
	.mem_to_bs_27 (mem_to_bs_27),
	.mem_to_bs_28 (mem_to_bs_28),
	.mem_to_bs_29 (mem_to_bs_29),
	.mem_to_bs_30 (mem_to_bs_30),
	.mem_to_bs_31 (mem_to_bs_31),
	.mem_to_bs_32 (mem_to_bs_32),
	.mem_to_bs_33 (mem_to_bs_33),
	.mem_to_bs_34 (mem_to_bs_34),
	.mem_to_bs_35 (mem_to_bs_35),
	.mem_to_bs_36 (mem_to_bs_36),
	.mem_to_bs_37 (mem_to_bs_37),
	.mem_to_bs_38 (mem_to_bs_38),
	.mem_to_bs_39 (mem_to_bs_39),
	.mem_to_bs_40 (mem_to_bs_40),
	.mem_to_bs_41 (mem_to_bs_41),
	.mem_to_bs_42 (mem_to_bs_42),
	.mem_to_bs_43 (mem_to_bs_43),
	.mem_to_bs_44 (mem_to_bs_44),
	.mem_to_bs_45 (mem_to_bs_45),
	.mem_to_bs_46 (mem_to_bs_46),
	.mem_to_bs_47 (mem_to_bs_47),
	.mem_to_bs_48 (mem_to_bs_48),
	.mem_to_bs_49 (mem_to_bs_49),
	.mem_to_bs_50 (mem_to_bs_50),
	.mem_to_bs_51 (mem_to_bs_51),
	.mem_to_bs_52 (mem_to_bs_52),
	.mem_to_bs_53 (mem_to_bs_53),
	.mem_to_bs_54 (mem_to_bs_54),
	.mem_to_bs_55 (mem_to_bs_55),
	.mem_to_bs_56 (mem_to_bs_56),
	.mem_to_bs_57 (mem_to_bs_57),
	.mem_to_bs_58 (mem_to_bs_58),
	.mem_to_bs_59 (mem_to_bs_59),
	.mem_to_bs_60 (mem_to_bs_60),
	.mem_to_bs_61 (mem_to_bs_61),
	.mem_to_bs_62 (mem_to_bs_62),
	.mem_to_bs_63 (mem_to_bs_63),
	.mem_to_bs_64 (mem_to_bs_64),
	.mem_to_bs_65 (mem_to_bs_65),
	.mem_to_bs_66 (mem_to_bs_66),
	.mem_to_bs_67 (mem_to_bs_67),
	.mem_to_bs_68 (mem_to_bs_68),
	.mem_to_bs_69 (mem_to_bs_69),
	.mem_to_bs_70 (mem_to_bs_70),
	.mem_to_bs_71 (mem_to_bs_71),
	.mem_to_bs_72 (mem_to_bs_72),
	.mem_to_bs_73 (mem_to_bs_73),
	.mem_to_bs_74 (mem_to_bs_74),
	.mem_to_bs_75 (mem_to_bs_75),
	.mem_to_bs_76 (mem_to_bs_76),
	.mem_to_bs_77 (mem_to_bs_77),
	.mem_to_bs_78 (mem_to_bs_78),
	.mem_to_bs_79 (mem_to_bs_79),
	.mem_to_bs_80 (mem_to_bs_80),
	.mem_to_bs_81 (mem_to_bs_81),
	.mem_to_bs_82 (mem_to_bs_82),
	.mem_to_bs_83 (mem_to_bs_83),
	.mem_to_bs_84 (mem_to_bs_84),
	// The memory Dout port to check nodes as instrinsic messages
	.mem_to_cnu_0  (mem_to_cnu_0 ),
	.mem_to_cnu_1  (mem_to_cnu_1 ),
	.mem_to_cnu_2  (mem_to_cnu_2 ),
	.mem_to_cnu_3  (mem_to_cnu_3 ),
	.mem_to_cnu_4  (mem_to_cnu_4 ),
	.mem_to_cnu_5  (mem_to_cnu_5 ),
	.mem_to_cnu_6  (mem_to_cnu_6 ),
	.mem_to_cnu_7  (mem_to_cnu_7 ),
	.mem_to_cnu_8  (mem_to_cnu_8 ),
	.mem_to_cnu_9  (mem_to_cnu_9 ),
	.mem_to_cnu_10 (mem_to_cnu_10),
	.mem_to_cnu_11 (mem_to_cnu_11),
	.mem_to_cnu_12 (mem_to_cnu_12),
	.mem_to_cnu_13 (mem_to_cnu_13),
	.mem_to_cnu_14 (mem_to_cnu_14),
	.mem_to_cnu_15 (mem_to_cnu_15),
	.mem_to_cnu_16 (mem_to_cnu_16),
	.mem_to_cnu_17 (mem_to_cnu_17),
	.mem_to_cnu_18 (mem_to_cnu_18),
	.mem_to_cnu_19 (mem_to_cnu_19),
	.mem_to_cnu_20 (mem_to_cnu_20),
	.mem_to_cnu_21 (mem_to_cnu_21),
	.mem_to_cnu_22 (mem_to_cnu_22),
	.mem_to_cnu_23 (mem_to_cnu_23),
	.mem_to_cnu_24 (mem_to_cnu_24),
	.mem_to_cnu_25 (mem_to_cnu_25),
	.mem_to_cnu_26 (mem_to_cnu_26),
	.mem_to_cnu_27 (mem_to_cnu_27),
	.mem_to_cnu_28 (mem_to_cnu_28),
	.mem_to_cnu_29 (mem_to_cnu_29),
	.mem_to_cnu_30 (mem_to_cnu_30),
	.mem_to_cnu_31 (mem_to_cnu_31),
	.mem_to_cnu_32 (mem_to_cnu_32),
	.mem_to_cnu_33 (mem_to_cnu_33),
	.mem_to_cnu_34 (mem_to_cnu_34),
	.mem_to_cnu_35 (mem_to_cnu_35),
	.mem_to_cnu_36 (mem_to_cnu_36),
	.mem_to_cnu_37 (mem_to_cnu_37),
	.mem_to_cnu_38 (mem_to_cnu_38),
	.mem_to_cnu_39 (mem_to_cnu_39),
	.mem_to_cnu_40 (mem_to_cnu_40),
	.mem_to_cnu_41 (mem_to_cnu_41),
	.mem_to_cnu_42 (mem_to_cnu_42),
	.mem_to_cnu_43 (mem_to_cnu_43),
	.mem_to_cnu_44 (mem_to_cnu_44),
	.mem_to_cnu_45 (mem_to_cnu_45),
	.mem_to_cnu_46 (mem_to_cnu_46),
	.mem_to_cnu_47 (mem_to_cnu_47),
	.mem_to_cnu_48 (mem_to_cnu_48),
	.mem_to_cnu_49 (mem_to_cnu_49),
	.mem_to_cnu_50 (mem_to_cnu_50),
	.mem_to_cnu_51 (mem_to_cnu_51),
	.mem_to_cnu_52 (mem_to_cnu_52),
	.mem_to_cnu_53 (mem_to_cnu_53),
	.mem_to_cnu_54 (mem_to_cnu_54),
	.mem_to_cnu_55 (mem_to_cnu_55),
	.mem_to_cnu_56 (mem_to_cnu_56),
	.mem_to_cnu_57 (mem_to_cnu_57),
	.mem_to_cnu_58 (mem_to_cnu_58),
	.mem_to_cnu_59 (mem_to_cnu_59),
	.mem_to_cnu_60 (mem_to_cnu_60),
	.mem_to_cnu_61 (mem_to_cnu_61),
	.mem_to_cnu_62 (mem_to_cnu_62),
	.mem_to_cnu_63 (mem_to_cnu_63),
	.mem_to_cnu_64 (mem_to_cnu_64),
	.mem_to_cnu_65 (mem_to_cnu_65),
	.mem_to_cnu_66 (mem_to_cnu_66),
	.mem_to_cnu_67 (mem_to_cnu_67),
	.mem_to_cnu_68 (mem_to_cnu_68),
	.mem_to_cnu_69 (mem_to_cnu_69),
	.mem_to_cnu_70 (mem_to_cnu_70),
	.mem_to_cnu_71 (mem_to_cnu_71),
	.mem_to_cnu_72 (mem_to_cnu_72),
	.mem_to_cnu_73 (mem_to_cnu_73),
	.mem_to_cnu_74 (mem_to_cnu_74),
	.mem_to_cnu_75 (mem_to_cnu_75),
	.mem_to_cnu_76 (mem_to_cnu_76),
	.mem_to_cnu_77 (mem_to_cnu_77),
	.mem_to_cnu_78 (mem_to_cnu_78),
	.mem_to_cnu_79 (mem_to_cnu_79),
	.mem_to_cnu_80 (mem_to_cnu_80),
	.mem_to_cnu_81 (mem_to_cnu_81),
	.mem_to_cnu_82 (mem_to_cnu_82),
	.mem_to_cnu_83 (mem_to_cnu_83),
	.mem_to_cnu_84 (mem_to_cnu_84),
	// From Dout port of extrinsic message RAMs
	.Din_0  (ram_dout_reg[0 ]),
	.Din_1  (ram_dout_reg[1 ]),
	.Din_2  (ram_dout_reg[2 ]),
	.Din_3  (ram_dout_reg[3 ]),
	.Din_4  (ram_dout_reg[4 ]),
	.Din_5  (ram_dout_reg[5 ]),
	.Din_6  (ram_dout_reg[6 ]),
	.Din_7  (ram_dout_reg[7 ]),
	.Din_8  (ram_dout_reg[8 ]),
	.Din_9  (ram_dout_reg[9 ]),
	.Din_10 (ram_dout_reg[10]),
	.Din_11 (ram_dout_reg[11]),
	.Din_12 (ram_dout_reg[12]),
	.Din_13 (ram_dout_reg[13]),
	.Din_14 (ram_dout_reg[14]),
	.Din_15 (ram_dout_reg[15]),
	.Din_16 (ram_dout_reg[16]),
	.Din_17 (ram_dout_reg[17]),
	.Din_18 (ram_dout_reg[18]),
	.Din_19 (ram_dout_reg[19]),
	.Din_20 (ram_dout_reg[20]),
	.Din_21 (ram_dout_reg[21]),
	.Din_22 (ram_dout_reg[22]),
	.Din_23 (ram_dout_reg[23]),
	.Din_24 (ram_dout_reg[24]),
	.Din_25 (ram_dout_reg[25]),
	.Din_26 (ram_dout_reg[26]),
	.Din_27 (ram_dout_reg[27]),
	.Din_28 (ram_dout_reg[28]),
	.Din_29 (ram_dout_reg[29]),
	.Din_30 (ram_dout_reg[30]),
	.Din_31 (ram_dout_reg[31]),
	.Din_32 (ram_dout_reg[32]),
	.Din_33 (ram_dout_reg[33]),
	.Din_34 (ram_dout_reg[34]),
	.Din_35 (ram_dout_reg[35]),
	.Din_36 (ram_dout_reg[36]),
	.Din_37 (ram_dout_reg[37]),
	.Din_38 (ram_dout_reg[38]),
	.Din_39 (ram_dout_reg[39]),
	.Din_40 (ram_dout_reg[40]),
	.Din_41 (ram_dout_reg[41]),
	.Din_42 (ram_dout_reg[42]),
	.Din_43 (ram_dout_reg[43]),
	.Din_44 (ram_dout_reg[44]),
	.Din_45 (ram_dout_reg[45]),
	.Din_46 (ram_dout_reg[46]),
	.Din_47 (ram_dout_reg[47]),
	.Din_48 (ram_dout_reg[48]),
	.Din_49 (ram_dout_reg[49]),
	.Din_50 (ram_dout_reg[50]),
	.Din_51 (ram_dout_reg[51]),
	.Din_52 (ram_dout_reg[52]),
	.Din_53 (ram_dout_reg[53]),
	.Din_54 (ram_dout_reg[54]),
	.Din_55 (ram_dout_reg[55]),
	.Din_56 (ram_dout_reg[56]),
	.Din_57 (ram_dout_reg[57]),
	.Din_58 (ram_dout_reg[58]),
	.Din_59 (ram_dout_reg[59]),
	.Din_60 (ram_dout_reg[60]),
	.Din_61 (ram_dout_reg[61]),
	.Din_62 (ram_dout_reg[62]),
	.Din_63 (ram_dout_reg[63]),
	.Din_64 (ram_dout_reg[64]),
	.Din_65 (ram_dout_reg[65]),
	.Din_66 (ram_dout_reg[66]),
	.Din_67 (ram_dout_reg[67]),
	.Din_68 (ram_dout_reg[68]),
	.Din_69 (ram_dout_reg[69]),
	.Din_70 (ram_dout_reg[70]),
	.Din_71 (ram_dout_reg[71]),
	.Din_72 (ram_dout_reg[72]),
	.Din_73 (ram_dout_reg[73]),
	.Din_74 (ram_dout_reg[74]),
	.Din_75 (ram_dout_reg[75]),
	.Din_76 (ram_dout_reg[76]),
	.Din_77 (ram_dout_reg[77]),
	.Din_78 (ram_dout_reg[78]),
	.Din_79 (ram_dout_reg[79]),
	.Din_80 (ram_dout_reg[80]),
	.Din_81 (ram_dout_reg[81]),
	.Din_82 (ram_dout_reg[82]),
	.Din_83 (ram_dout_reg[83]),
	.Din_84 (ram_dout_reg[84]),

	.sched_cmd (sched_cmd) // 1'b0: align_in from variable msg; 1'b1: align_in from check msg
);
endmodule

module ram_out_demux #(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 85
) (
	// The memory Dout port to permutation network for instrinsic messages of variable nodes of upcoming operation
	output wire [QUAN_SIZE-1:0] mem_to_bs_0,
	output wire [QUAN_SIZE-1:0] mem_to_bs_1,
	output wire [QUAN_SIZE-1:0] mem_to_bs_2,
	output wire [QUAN_SIZE-1:0] mem_to_bs_3,
	output wire [QUAN_SIZE-1:0] mem_to_bs_4,
	output wire [QUAN_SIZE-1:0] mem_to_bs_5,
	output wire [QUAN_SIZE-1:0] mem_to_bs_6,
	output wire [QUAN_SIZE-1:0] mem_to_bs_7,
	output wire [QUAN_SIZE-1:0] mem_to_bs_8,
	output wire [QUAN_SIZE-1:0] mem_to_bs_9,
	output wire [QUAN_SIZE-1:0] mem_to_bs_10,
	output wire [QUAN_SIZE-1:0] mem_to_bs_11,
	output wire [QUAN_SIZE-1:0] mem_to_bs_12,
	output wire [QUAN_SIZE-1:0] mem_to_bs_13,
	output wire [QUAN_SIZE-1:0] mem_to_bs_14,
	output wire [QUAN_SIZE-1:0] mem_to_bs_15,
	output wire [QUAN_SIZE-1:0] mem_to_bs_16,
	output wire [QUAN_SIZE-1:0] mem_to_bs_17,
	output wire [QUAN_SIZE-1:0] mem_to_bs_18,
	output wire [QUAN_SIZE-1:0] mem_to_bs_19,
	output wire [QUAN_SIZE-1:0] mem_to_bs_20,
	output wire [QUAN_SIZE-1:0] mem_to_bs_21,
	output wire [QUAN_SIZE-1:0] mem_to_bs_22,
	output wire [QUAN_SIZE-1:0] mem_to_bs_23,
	output wire [QUAN_SIZE-1:0] mem_to_bs_24,
	output wire [QUAN_SIZE-1:0] mem_to_bs_25,
	output wire [QUAN_SIZE-1:0] mem_to_bs_26,
	output wire [QUAN_SIZE-1:0] mem_to_bs_27,
	output wire [QUAN_SIZE-1:0] mem_to_bs_28,
	output wire [QUAN_SIZE-1:0] mem_to_bs_29,
	output wire [QUAN_SIZE-1:0] mem_to_bs_30,
	output wire [QUAN_SIZE-1:0] mem_to_bs_31,
	output wire [QUAN_SIZE-1:0] mem_to_bs_32,
	output wire [QUAN_SIZE-1:0] mem_to_bs_33,
	output wire [QUAN_SIZE-1:0] mem_to_bs_34,
	output wire [QUAN_SIZE-1:0] mem_to_bs_35,
	output wire [QUAN_SIZE-1:0] mem_to_bs_36,
	output wire [QUAN_SIZE-1:0] mem_to_bs_37,
	output wire [QUAN_SIZE-1:0] mem_to_bs_38,
	output wire [QUAN_SIZE-1:0] mem_to_bs_39,
	output wire [QUAN_SIZE-1:0] mem_to_bs_40,
	output wire [QUAN_SIZE-1:0] mem_to_bs_41,
	output wire [QUAN_SIZE-1:0] mem_to_bs_42,
	output wire [QUAN_SIZE-1:0] mem_to_bs_43,
	output wire [QUAN_SIZE-1:0] mem_to_bs_44,
	output wire [QUAN_SIZE-1:0] mem_to_bs_45,
	output wire [QUAN_SIZE-1:0] mem_to_bs_46,
	output wire [QUAN_SIZE-1:0] mem_to_bs_47,
	output wire [QUAN_SIZE-1:0] mem_to_bs_48,
	output wire [QUAN_SIZE-1:0] mem_to_bs_49,
	output wire [QUAN_SIZE-1:0] mem_to_bs_50,
	output wire [QUAN_SIZE-1:0] mem_to_bs_51,
	output wire [QUAN_SIZE-1:0] mem_to_bs_52,
	output wire [QUAN_SIZE-1:0] mem_to_bs_53,
	output wire [QUAN_SIZE-1:0] mem_to_bs_54,
	output wire [QUAN_SIZE-1:0] mem_to_bs_55,
	output wire [QUAN_SIZE-1:0] mem_to_bs_56,
	output wire [QUAN_SIZE-1:0] mem_to_bs_57,
	output wire [QUAN_SIZE-1:0] mem_to_bs_58,
	output wire [QUAN_SIZE-1:0] mem_to_bs_59,
	output wire [QUAN_SIZE-1:0] mem_to_bs_60,
	output wire [QUAN_SIZE-1:0] mem_to_bs_61,
	output wire [QUAN_SIZE-1:0] mem_to_bs_62,
	output wire [QUAN_SIZE-1:0] mem_to_bs_63,
	output wire [QUAN_SIZE-1:0] mem_to_bs_64,
	output wire [QUAN_SIZE-1:0] mem_to_bs_65,
	output wire [QUAN_SIZE-1:0] mem_to_bs_66,
	output wire [QUAN_SIZE-1:0] mem_to_bs_67,
	output wire [QUAN_SIZE-1:0] mem_to_bs_68,
	output wire [QUAN_SIZE-1:0] mem_to_bs_69,
	output wire [QUAN_SIZE-1:0] mem_to_bs_70,
	output wire [QUAN_SIZE-1:0] mem_to_bs_71,
	output wire [QUAN_SIZE-1:0] mem_to_bs_72,
	output wire [QUAN_SIZE-1:0] mem_to_bs_73,
	output wire [QUAN_SIZE-1:0] mem_to_bs_74,
	output wire [QUAN_SIZE-1:0] mem_to_bs_75,
	output wire [QUAN_SIZE-1:0] mem_to_bs_76,
	output wire [QUAN_SIZE-1:0] mem_to_bs_77,
	output wire [QUAN_SIZE-1:0] mem_to_bs_78,
	output wire [QUAN_SIZE-1:0] mem_to_bs_79,
	output wire [QUAN_SIZE-1:0] mem_to_bs_80,
	output wire [QUAN_SIZE-1:0] mem_to_bs_81,
	output wire [QUAN_SIZE-1:0] mem_to_bs_82,
	output wire [QUAN_SIZE-1:0] mem_to_bs_83,
	output wire [QUAN_SIZE-1:0] mem_to_bs_84,
	// The memory Dout port to check nodes as instrinsic messages
	output wire [QUAN_SIZE-1:0] mem_to_cnu_0,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_1,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_2,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_3,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_4,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_5,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_6,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_7,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_8,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_9,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_10,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_11,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_12,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_13,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_14,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_15,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_16,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_17,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_18,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_19,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_20,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_21,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_22,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_23,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_24,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_25,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_26,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_27,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_28,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_29,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_30,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_31,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_32,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_33,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_34,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_35,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_36,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_37,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_38,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_39,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_40,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_41,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_42,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_43,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_44,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_45,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_46,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_47,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_48,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_49,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_50,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_51,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_52,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_53,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_54,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_55,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_56,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_57,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_58,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_59,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_60,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_61,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_62,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_63,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_64,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_65,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_66,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_67,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_68,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_69,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_70,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_71,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_72,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_73,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_74,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_75,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_76,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_77,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_78,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_79,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_80,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_81,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_82,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_83,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_84,
	// From Dout port of extrinsic message RAMs
	input wire [QUAN_SIZE-1:0] Din_0,
	input wire [QUAN_SIZE-1:0] Din_1,
	input wire [QUAN_SIZE-1:0] Din_2,
	input wire [QUAN_SIZE-1:0] Din_3,
	input wire [QUAN_SIZE-1:0] Din_4,
	input wire [QUAN_SIZE-1:0] Din_5,
	input wire [QUAN_SIZE-1:0] Din_6,
	input wire [QUAN_SIZE-1:0] Din_7,
	input wire [QUAN_SIZE-1:0] Din_8,
	input wire [QUAN_SIZE-1:0] Din_9,
	input wire [QUAN_SIZE-1:0] Din_10,
	input wire [QUAN_SIZE-1:0] Din_11,
	input wire [QUAN_SIZE-1:0] Din_12,
	input wire [QUAN_SIZE-1:0] Din_13,
	input wire [QUAN_SIZE-1:0] Din_14,
	input wire [QUAN_SIZE-1:0] Din_15,
	input wire [QUAN_SIZE-1:0] Din_16,
	input wire [QUAN_SIZE-1:0] Din_17,
	input wire [QUAN_SIZE-1:0] Din_18,
	input wire [QUAN_SIZE-1:0] Din_19,
	input wire [QUAN_SIZE-1:0] Din_20,
	input wire [QUAN_SIZE-1:0] Din_21,
	input wire [QUAN_SIZE-1:0] Din_22,
	input wire [QUAN_SIZE-1:0] Din_23,
	input wire [QUAN_SIZE-1:0] Din_24,
	input wire [QUAN_SIZE-1:0] Din_25,
	input wire [QUAN_SIZE-1:0] Din_26,
	input wire [QUAN_SIZE-1:0] Din_27,
	input wire [QUAN_SIZE-1:0] Din_28,
	input wire [QUAN_SIZE-1:0] Din_29,
	input wire [QUAN_SIZE-1:0] Din_30,
	input wire [QUAN_SIZE-1:0] Din_31,
	input wire [QUAN_SIZE-1:0] Din_32,
	input wire [QUAN_SIZE-1:0] Din_33,
	input wire [QUAN_SIZE-1:0] Din_34,
	input wire [QUAN_SIZE-1:0] Din_35,
	input wire [QUAN_SIZE-1:0] Din_36,
	input wire [QUAN_SIZE-1:0] Din_37,
	input wire [QUAN_SIZE-1:0] Din_38,
	input wire [QUAN_SIZE-1:0] Din_39,
	input wire [QUAN_SIZE-1:0] Din_40,
	input wire [QUAN_SIZE-1:0] Din_41,
	input wire [QUAN_SIZE-1:0] Din_42,
	input wire [QUAN_SIZE-1:0] Din_43,
	input wire [QUAN_SIZE-1:0] Din_44,
	input wire [QUAN_SIZE-1:0] Din_45,
	input wire [QUAN_SIZE-1:0] Din_46,
	input wire [QUAN_SIZE-1:0] Din_47,
	input wire [QUAN_SIZE-1:0] Din_48,
	input wire [QUAN_SIZE-1:0] Din_49,
	input wire [QUAN_SIZE-1:0] Din_50,
	input wire [QUAN_SIZE-1:0] Din_51,
	input wire [QUAN_SIZE-1:0] Din_52,
	input wire [QUAN_SIZE-1:0] Din_53,
	input wire [QUAN_SIZE-1:0] Din_54,
	input wire [QUAN_SIZE-1:0] Din_55,
	input wire [QUAN_SIZE-1:0] Din_56,
	input wire [QUAN_SIZE-1:0] Din_57,
	input wire [QUAN_SIZE-1:0] Din_58,
	input wire [QUAN_SIZE-1:0] Din_59,
	input wire [QUAN_SIZE-1:0] Din_60,
	input wire [QUAN_SIZE-1:0] Din_61,
	input wire [QUAN_SIZE-1:0] Din_62,
	input wire [QUAN_SIZE-1:0] Din_63,
	input wire [QUAN_SIZE-1:0] Din_64,
	input wire [QUAN_SIZE-1:0] Din_65,
	input wire [QUAN_SIZE-1:0] Din_66,
	input wire [QUAN_SIZE-1:0] Din_67,
	input wire [QUAN_SIZE-1:0] Din_68,
	input wire [QUAN_SIZE-1:0] Din_69,
	input wire [QUAN_SIZE-1:0] Din_70,
	input wire [QUAN_SIZE-1:0] Din_71,
	input wire [QUAN_SIZE-1:0] Din_72,
	input wire [QUAN_SIZE-1:0] Din_73,
	input wire [QUAN_SIZE-1:0] Din_74,
	input wire [QUAN_SIZE-1:0] Din_75,
	input wire [QUAN_SIZE-1:0] Din_76,
	input wire [QUAN_SIZE-1:0] Din_77,
	input wire [QUAN_SIZE-1:0] Din_78,
	input wire [QUAN_SIZE-1:0] Din_79,
	input wire [QUAN_SIZE-1:0] Din_80,
	input wire [QUAN_SIZE-1:0] Din_81,
	input wire [QUAN_SIZE-1:0] Din_82,
	input wire [QUAN_SIZE-1:0] Din_83,
	input wire [QUAN_SIZE-1:0] Din_84,

	input wire sched_cmd // 1'b0: align_in from variable msg; 1'b1: align_in from check msg
);

assign mem_to_bs_0 = (sched_cmd == 1'b1) ? Din_0 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_1 = (sched_cmd == 1'b1) ? Din_1 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_2 = (sched_cmd == 1'b1) ? Din_2 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_3 = (sched_cmd == 1'b1) ? Din_3 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_4 = (sched_cmd == 1'b1) ? Din_4 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_5 = (sched_cmd == 1'b1) ? Din_5 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_6 = (sched_cmd == 1'b1) ? Din_6 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_7 = (sched_cmd == 1'b1) ? Din_7 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_8 = (sched_cmd == 1'b1) ? Din_8 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_9 = (sched_cmd == 1'b1) ? Din_9 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_10 = (sched_cmd == 1'b1) ? Din_10 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_11 = (sched_cmd == 1'b1) ? Din_11 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_12 = (sched_cmd == 1'b1) ? Din_12 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_13 = (sched_cmd == 1'b1) ? Din_13 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_14 = (sched_cmd == 1'b1) ? Din_14 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_15 = (sched_cmd == 1'b1) ? Din_15 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_16 = (sched_cmd == 1'b1) ? Din_16 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_17 = (sched_cmd == 1'b1) ? Din_17 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_18 = (sched_cmd == 1'b1) ? Din_18 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_19 = (sched_cmd == 1'b1) ? Din_19 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_20 = (sched_cmd == 1'b1) ? Din_20 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_21 = (sched_cmd == 1'b1) ? Din_21 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_22 = (sched_cmd == 1'b1) ? Din_22 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_23 = (sched_cmd == 1'b1) ? Din_23 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_24 = (sched_cmd == 1'b1) ? Din_24 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_25 = (sched_cmd == 1'b1) ? Din_25 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_26 = (sched_cmd == 1'b1) ? Din_26 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_27 = (sched_cmd == 1'b1) ? Din_27 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_28 = (sched_cmd == 1'b1) ? Din_28 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_29 = (sched_cmd == 1'b1) ? Din_29 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_30 = (sched_cmd == 1'b1) ? Din_30 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_31 = (sched_cmd == 1'b1) ? Din_31 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_32 = (sched_cmd == 1'b1) ? Din_32 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_33 = (sched_cmd == 1'b1) ? Din_33 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_34 = (sched_cmd == 1'b1) ? Din_34 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_35 = (sched_cmd == 1'b1) ? Din_35 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_36 = (sched_cmd == 1'b1) ? Din_36 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_37 = (sched_cmd == 1'b1) ? Din_37 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_38 = (sched_cmd == 1'b1) ? Din_38 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_39 = (sched_cmd == 1'b1) ? Din_39 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_40 = (sched_cmd == 1'b1) ? Din_40 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_41 = (sched_cmd == 1'b1) ? Din_41 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_42 = (sched_cmd == 1'b1) ? Din_42 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_43 = (sched_cmd == 1'b1) ? Din_43 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_44 = (sched_cmd == 1'b1) ? Din_44 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_45 = (sched_cmd == 1'b1) ? Din_45 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_46 = (sched_cmd == 1'b1) ? Din_46 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_47 = (sched_cmd == 1'b1) ? Din_47 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_48 = (sched_cmd == 1'b1) ? Din_48 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_49 = (sched_cmd == 1'b1) ? Din_49 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_50 = (sched_cmd == 1'b1) ? Din_50 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_51 = (sched_cmd == 1'b1) ? Din_51 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_52 = (sched_cmd == 1'b1) ? Din_52 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_53 = (sched_cmd == 1'b1) ? Din_53 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_54 = (sched_cmd == 1'b1) ? Din_54 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_55 = (sched_cmd == 1'b1) ? Din_55 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_56 = (sched_cmd == 1'b1) ? Din_56 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_57 = (sched_cmd == 1'b1) ? Din_57 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_58 = (sched_cmd == 1'b1) ? Din_58 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_59 = (sched_cmd == 1'b1) ? Din_59 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_60 = (sched_cmd == 1'b1) ? Din_60 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_61 = (sched_cmd == 1'b1) ? Din_61 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_62 = (sched_cmd == 1'b1) ? Din_62 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_63 = (sched_cmd == 1'b1) ? Din_63 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_64 = (sched_cmd == 1'b1) ? Din_64 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_65 = (sched_cmd == 1'b1) ? Din_65 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_66 = (sched_cmd == 1'b1) ? Din_66 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_67 = (sched_cmd == 1'b1) ? Din_67 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_68 = (sched_cmd == 1'b1) ? Din_68 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_69 = (sched_cmd == 1'b1) ? Din_69 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_70 = (sched_cmd == 1'b1) ? Din_70 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_71 = (sched_cmd == 1'b1) ? Din_71 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_72 = (sched_cmd == 1'b1) ? Din_72 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_73 = (sched_cmd == 1'b1) ? Din_73 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_74 = (sched_cmd == 1'b1) ? Din_74 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_75 = (sched_cmd == 1'b1) ? Din_75 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_76 = (sched_cmd == 1'b1) ? Din_76 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_77 = (sched_cmd == 1'b1) ? Din_77 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_78 = (sched_cmd == 1'b1) ? Din_78 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_79 = (sched_cmd == 1'b1) ? Din_79 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_80 = (sched_cmd == 1'b1) ? Din_80 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_81 = (sched_cmd == 1'b1) ? Din_81 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_82 = (sched_cmd == 1'b1) ? Din_82 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_83 = (sched_cmd == 1'b1) ? Din_83 : {QUAN_SIZE{1'bz}};
assign mem_to_bs_84 = (sched_cmd == 1'b1) ? Din_84 : {QUAN_SIZE{1'bz}};

assign mem_to_cnu_0 = (sched_cmd == 1'b0) ? Din_0 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_1 = (sched_cmd == 1'b0) ? Din_1 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_2 = (sched_cmd == 1'b0) ? Din_2 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_3 = (sched_cmd == 1'b0) ? Din_3 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_4 = (sched_cmd == 1'b0) ? Din_4 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_5 = (sched_cmd == 1'b0) ? Din_5 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_6 = (sched_cmd == 1'b0) ? Din_6 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_7 = (sched_cmd == 1'b0) ? Din_7 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_8 = (sched_cmd == 1'b0) ? Din_8 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_9 = (sched_cmd == 1'b0) ? Din_9 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_10 = (sched_cmd == 1'b0) ? Din_10 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_11 = (sched_cmd == 1'b0) ? Din_11 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_12 = (sched_cmd == 1'b0) ? Din_12 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_13 = (sched_cmd == 1'b0) ? Din_13 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_14 = (sched_cmd == 1'b0) ? Din_14 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_15 = (sched_cmd == 1'b0) ? Din_15 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_16 = (sched_cmd == 1'b0) ? Din_16 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_17 = (sched_cmd == 1'b0) ? Din_17 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_18 = (sched_cmd == 1'b0) ? Din_18 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_19 = (sched_cmd == 1'b0) ? Din_19 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_20 = (sched_cmd == 1'b0) ? Din_20 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_21 = (sched_cmd == 1'b0) ? Din_21 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_22 = (sched_cmd == 1'b0) ? Din_22 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_23 = (sched_cmd == 1'b0) ? Din_23 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_24 = (sched_cmd == 1'b0) ? Din_24 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_25 = (sched_cmd == 1'b0) ? Din_25 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_26 = (sched_cmd == 1'b0) ? Din_26 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_27 = (sched_cmd == 1'b0) ? Din_27 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_28 = (sched_cmd == 1'b0) ? Din_28 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_29 = (sched_cmd == 1'b0) ? Din_29 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_30 = (sched_cmd == 1'b0) ? Din_30 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_31 = (sched_cmd == 1'b0) ? Din_31 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_32 = (sched_cmd == 1'b0) ? Din_32 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_33 = (sched_cmd == 1'b0) ? Din_33 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_34 = (sched_cmd == 1'b0) ? Din_34 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_35 = (sched_cmd == 1'b0) ? Din_35 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_36 = (sched_cmd == 1'b0) ? Din_36 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_37 = (sched_cmd == 1'b0) ? Din_37 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_38 = (sched_cmd == 1'b0) ? Din_38 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_39 = (sched_cmd == 1'b0) ? Din_39 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_40 = (sched_cmd == 1'b0) ? Din_40 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_41 = (sched_cmd == 1'b0) ? Din_41 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_42 = (sched_cmd == 1'b0) ? Din_42 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_43 = (sched_cmd == 1'b0) ? Din_43 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_44 = (sched_cmd == 1'b0) ? Din_44 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_45 = (sched_cmd == 1'b0) ? Din_45 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_46 = (sched_cmd == 1'b0) ? Din_46 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_47 = (sched_cmd == 1'b0) ? Din_47 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_48 = (sched_cmd == 1'b0) ? Din_48 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_49 = (sched_cmd == 1'b0) ? Din_49 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_50 = (sched_cmd == 1'b0) ? Din_50 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_51 = (sched_cmd == 1'b0) ? Din_51 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_52 = (sched_cmd == 1'b0) ? Din_52 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_53 = (sched_cmd == 1'b0) ? Din_53 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_54 = (sched_cmd == 1'b0) ? Din_54 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_55 = (sched_cmd == 1'b0) ? Din_55 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_56 = (sched_cmd == 1'b0) ? Din_56 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_57 = (sched_cmd == 1'b0) ? Din_57 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_58 = (sched_cmd == 1'b0) ? Din_58 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_59 = (sched_cmd == 1'b0) ? Din_59 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_60 = (sched_cmd == 1'b0) ? Din_60 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_61 = (sched_cmd == 1'b0) ? Din_61 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_62 = (sched_cmd == 1'b0) ? Din_62 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_63 = (sched_cmd == 1'b0) ? Din_63 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_64 = (sched_cmd == 1'b0) ? Din_64 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_65 = (sched_cmd == 1'b0) ? Din_65 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_66 = (sched_cmd == 1'b0) ? Din_66 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_67 = (sched_cmd == 1'b0) ? Din_67 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_68 = (sched_cmd == 1'b0) ? Din_68 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_69 = (sched_cmd == 1'b0) ? Din_69 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_70 = (sched_cmd == 1'b0) ? Din_70 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_71 = (sched_cmd == 1'b0) ? Din_71 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_72 = (sched_cmd == 1'b0) ? Din_72 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_73 = (sched_cmd == 1'b0) ? Din_73 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_74 = (sched_cmd == 1'b0) ? Din_74 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_75 = (sched_cmd == 1'b0) ? Din_75 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_76 = (sched_cmd == 1'b0) ? Din_76 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_77 = (sched_cmd == 1'b0) ? Din_77 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_78 = (sched_cmd == 1'b0) ? Din_78 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_79 = (sched_cmd == 1'b0) ? Din_79 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_80 = (sched_cmd == 1'b0) ? Din_80 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_81 = (sched_cmd == 1'b0) ? Din_81 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_82 = (sched_cmd == 1'b0) ? Din_82 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_83 = (sched_cmd == 1'b0) ? Din_83 : {QUAN_SIZE{1'bz}};
assign mem_to_cnu_84 = (sched_cmd == 1'b0) ? Din_84 : {QUAN_SIZE{1'bz}};
endmodule