`include "define.vh"

`ifdef SCHED_4_6
module ram_pageAlign_interface_submatrix_0#(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 85,
	parameter LAYER_NUM = 3
) (
	output reg [QUAN_SIZE-1:0] msg_out_0,
	output reg [QUAN_SIZE-1:0] msg_out_1,
	output reg [QUAN_SIZE-1:0] msg_out_2,
	output reg [QUAN_SIZE-1:0] msg_out_3,
	output reg [QUAN_SIZE-1:0] msg_out_4,
	output reg [QUAN_SIZE-1:0] msg_out_5,
	output reg [QUAN_SIZE-1:0] msg_out_6,
	output reg [QUAN_SIZE-1:0] msg_out_7,
	output reg [QUAN_SIZE-1:0] msg_out_8,
	output reg [QUAN_SIZE-1:0] msg_out_9,
	output reg [QUAN_SIZE-1:0] msg_out_10,
	output reg [QUAN_SIZE-1:0] msg_out_11,
	output reg [QUAN_SIZE-1:0] msg_out_12,
	output reg [QUAN_SIZE-1:0] msg_out_13,
	output reg [QUAN_SIZE-1:0] msg_out_14,
	output reg [QUAN_SIZE-1:0] msg_out_15,
	output reg [QUAN_SIZE-1:0] msg_out_16,
	output reg [QUAN_SIZE-1:0] msg_out_17,
	output reg [QUAN_SIZE-1:0] msg_out_18,
	output reg [QUAN_SIZE-1:0] msg_out_19,
	output reg [QUAN_SIZE-1:0] msg_out_20,
	output reg [QUAN_SIZE-1:0] msg_out_21,
	output reg [QUAN_SIZE-1:0] msg_out_22,
	output reg [QUAN_SIZE-1:0] msg_out_23,
	output reg [QUAN_SIZE-1:0] msg_out_24,
	output reg [QUAN_SIZE-1:0] msg_out_25,
	output reg [QUAN_SIZE-1:0] msg_out_26,
	output reg [QUAN_SIZE-1:0] msg_out_27,
	output reg [QUAN_SIZE-1:0] msg_out_28,
	output reg [QUAN_SIZE-1:0] msg_out_29,
	output reg [QUAN_SIZE-1:0] msg_out_30,
	output reg [QUAN_SIZE-1:0] msg_out_31,
	output reg [QUAN_SIZE-1:0] msg_out_32,
	output reg [QUAN_SIZE-1:0] msg_out_33,
	output reg [QUAN_SIZE-1:0] msg_out_34,
	output reg [QUAN_SIZE-1:0] msg_out_35,
	output reg [QUAN_SIZE-1:0] msg_out_36,
	output reg [QUAN_SIZE-1:0] msg_out_37,
	output reg [QUAN_SIZE-1:0] msg_out_38,
	output reg [QUAN_SIZE-1:0] msg_out_39,
	output reg [QUAN_SIZE-1:0] msg_out_40,
	output reg [QUAN_SIZE-1:0] msg_out_41,
	output reg [QUAN_SIZE-1:0] msg_out_42,
	output reg [QUAN_SIZE-1:0] msg_out_43,
	output reg [QUAN_SIZE-1:0] msg_out_44,
	output reg [QUAN_SIZE-1:0] msg_out_45,
	output reg [QUAN_SIZE-1:0] msg_out_46,
	output reg [QUAN_SIZE-1:0] msg_out_47,
	output reg [QUAN_SIZE-1:0] msg_out_48,
	output reg [QUAN_SIZE-1:0] msg_out_49,
	output reg [QUAN_SIZE-1:0] msg_out_50,
	output reg [QUAN_SIZE-1:0] msg_out_51,
	output reg [QUAN_SIZE-1:0] msg_out_52,
	output reg [QUAN_SIZE-1:0] msg_out_53,
	output reg [QUAN_SIZE-1:0] msg_out_54,
	output reg [QUAN_SIZE-1:0] msg_out_55,
	output reg [QUAN_SIZE-1:0] msg_out_56,
	output reg [QUAN_SIZE-1:0] msg_out_57,
	output reg [QUAN_SIZE-1:0] msg_out_58,
	output reg [QUAN_SIZE-1:0] msg_out_59,
	output reg [QUAN_SIZE-1:0] msg_out_60,
	output reg [QUAN_SIZE-1:0] msg_out_61,
	output reg [QUAN_SIZE-1:0] msg_out_62,
	output reg [QUAN_SIZE-1:0] msg_out_63,
	output reg [QUAN_SIZE-1:0] msg_out_64,
	output reg [QUAN_SIZE-1:0] msg_out_65,
	output reg [QUAN_SIZE-1:0] msg_out_66,
	output reg [QUAN_SIZE-1:0] msg_out_67,
	output reg [QUAN_SIZE-1:0] msg_out_68,
	output reg [QUAN_SIZE-1:0] msg_out_69,
	output reg [QUAN_SIZE-1:0] msg_out_70,
	output reg [QUAN_SIZE-1:0] msg_out_71,
	output reg [QUAN_SIZE-1:0] msg_out_72,
	output reg [QUAN_SIZE-1:0] msg_out_73,
	output reg [QUAN_SIZE-1:0] msg_out_74,
	output reg [QUAN_SIZE-1:0] msg_out_75,
	output reg [QUAN_SIZE-1:0] msg_out_76,
	output reg [QUAN_SIZE-1:0] msg_out_77,
	output reg [QUAN_SIZE-1:0] msg_out_78,
	output reg [QUAN_SIZE-1:0] msg_out_79,
	output reg [QUAN_SIZE-1:0] msg_out_80,
	output reg [QUAN_SIZE-1:0] msg_out_81,
	output reg [QUAN_SIZE-1:0] msg_out_82,
	output reg [QUAN_SIZE-1:0] msg_out_83,
	output reg [QUAN_SIZE-1:0] msg_out_84,

	input wire [QUAN_SIZE-1:0] msg_in_0,
	input wire [QUAN_SIZE-1:0] msg_in_1,
	input wire [QUAN_SIZE-1:0] msg_in_2,
	input wire [QUAN_SIZE-1:0] msg_in_3,
	input wire [QUAN_SIZE-1:0] msg_in_4,
	input wire [QUAN_SIZE-1:0] msg_in_5,
	input wire [QUAN_SIZE-1:0] msg_in_6,
	input wire [QUAN_SIZE-1:0] msg_in_7,
	input wire [QUAN_SIZE-1:0] msg_in_8,
	input wire [QUAN_SIZE-1:0] msg_in_9,
	input wire [QUAN_SIZE-1:0] msg_in_10,
	input wire [QUAN_SIZE-1:0] msg_in_11,
	input wire [QUAN_SIZE-1:0] msg_in_12,
	input wire [QUAN_SIZE-1:0] msg_in_13,
	input wire [QUAN_SIZE-1:0] msg_in_14,
	input wire [QUAN_SIZE-1:0] msg_in_15,
	input wire [QUAN_SIZE-1:0] msg_in_16,
	input wire [QUAN_SIZE-1:0] msg_in_17,
	input wire [QUAN_SIZE-1:0] msg_in_18,
	input wire [QUAN_SIZE-1:0] msg_in_19,
	input wire [QUAN_SIZE-1:0] msg_in_20,
	input wire [QUAN_SIZE-1:0] msg_in_21,
	input wire [QUAN_SIZE-1:0] msg_in_22,
	input wire [QUAN_SIZE-1:0] msg_in_23,
	input wire [QUAN_SIZE-1:0] msg_in_24,
	input wire [QUAN_SIZE-1:0] msg_in_25,
	input wire [QUAN_SIZE-1:0] msg_in_26,
	input wire [QUAN_SIZE-1:0] msg_in_27,
	input wire [QUAN_SIZE-1:0] msg_in_28,
	input wire [QUAN_SIZE-1:0] msg_in_29,
	input wire [QUAN_SIZE-1:0] msg_in_30,
	input wire [QUAN_SIZE-1:0] msg_in_31,
	input wire [QUAN_SIZE-1:0] msg_in_32,
	input wire [QUAN_SIZE-1:0] msg_in_33,
	input wire [QUAN_SIZE-1:0] msg_in_34,
	input wire [QUAN_SIZE-1:0] msg_in_35,
	input wire [QUAN_SIZE-1:0] msg_in_36,
	input wire [QUAN_SIZE-1:0] msg_in_37,
	input wire [QUAN_SIZE-1:0] msg_in_38,
	input wire [QUAN_SIZE-1:0] msg_in_39,
	input wire [QUAN_SIZE-1:0] msg_in_40,
	input wire [QUAN_SIZE-1:0] msg_in_41,
	input wire [QUAN_SIZE-1:0] msg_in_42,
	input wire [QUAN_SIZE-1:0] msg_in_43,
	input wire [QUAN_SIZE-1:0] msg_in_44,
	input wire [QUAN_SIZE-1:0] msg_in_45,
	input wire [QUAN_SIZE-1:0] msg_in_46,
	input wire [QUAN_SIZE-1:0] msg_in_47,
	input wire [QUAN_SIZE-1:0] msg_in_48,
	input wire [QUAN_SIZE-1:0] msg_in_49,
	input wire [QUAN_SIZE-1:0] msg_in_50,
	input wire [QUAN_SIZE-1:0] msg_in_51,
	input wire [QUAN_SIZE-1:0] msg_in_52,
	input wire [QUAN_SIZE-1:0] msg_in_53,
	input wire [QUAN_SIZE-1:0] msg_in_54,
	input wire [QUAN_SIZE-1:0] msg_in_55,
	input wire [QUAN_SIZE-1:0] msg_in_56,
	input wire [QUAN_SIZE-1:0] msg_in_57,
	input wire [QUAN_SIZE-1:0] msg_in_58,
	input wire [QUAN_SIZE-1:0] msg_in_59,
	input wire [QUAN_SIZE-1:0] msg_in_60,
	input wire [QUAN_SIZE-1:0] msg_in_61,
	input wire [QUAN_SIZE-1:0] msg_in_62,
	input wire [QUAN_SIZE-1:0] msg_in_63,
	input wire [QUAN_SIZE-1:0] msg_in_64,
	input wire [QUAN_SIZE-1:0] msg_in_65,
	input wire [QUAN_SIZE-1:0] msg_in_66,
	input wire [QUAN_SIZE-1:0] msg_in_67,
	input wire [QUAN_SIZE-1:0] msg_in_68,
	input wire [QUAN_SIZE-1:0] msg_in_69,
	input wire [QUAN_SIZE-1:0] msg_in_70,
	input wire [QUAN_SIZE-1:0] msg_in_71,
	input wire [QUAN_SIZE-1:0] msg_in_72,
	input wire [QUAN_SIZE-1:0] msg_in_73,
	input wire [QUAN_SIZE-1:0] msg_in_74,
	input wire [QUAN_SIZE-1:0] msg_in_75,
	input wire [QUAN_SIZE-1:0] msg_in_76,
	input wire [QUAN_SIZE-1:0] msg_in_77,
	input wire [QUAN_SIZE-1:0] msg_in_78,
	input wire [QUAN_SIZE-1:0] msg_in_79,
	input wire [QUAN_SIZE-1:0] msg_in_80,
	input wire [QUAN_SIZE-1:0] msg_in_81,
	input wire [QUAN_SIZE-1:0] msg_in_82,
	input wire [QUAN_SIZE-1:0] msg_in_83,
	input wire [QUAN_SIZE-1:0] msg_in_84,

	input wire [LAYER_NUM-1:0] layer_status,
	input wire first_row_chunk,
	input wire sys_clk,
	input wire rstn
);

always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_0 <= 0; else msg_out_0 <= msg_in_0; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_1 <= 0; else msg_out_1 <= msg_in_1; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_2 <= 0; else msg_out_2 <= msg_in_2; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_3 <= 0; else msg_out_3 <= msg_in_3; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_4 <= 0; else msg_out_4 <= msg_in_4; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_5 <= 0; else msg_out_5 <= msg_in_5; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_6 <= 0; else msg_out_6 <= msg_in_6; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_7 <= 0; else msg_out_7 <= msg_in_7; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_8 <= 0; else msg_out_8 <= msg_in_8; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_9 <= 0; else msg_out_9 <= msg_in_9; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_10 <= 0; else msg_out_10 <= msg_in_10; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_11 <= 0; else msg_out_11 <= msg_in_11; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_12 <= 0; else msg_out_12 <= msg_in_12; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_13 <= 0; else msg_out_13 <= msg_in_13; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_14 <= 0; else msg_out_14 <= msg_in_14; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_15 <= 0; else msg_out_15 <= msg_in_15; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_16 <= 0; else msg_out_16 <= msg_in_16; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_17 <= 0; else msg_out_17 <= msg_in_17; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_18 <= 0; else msg_out_18 <= msg_in_18; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_19 <= 0; else msg_out_19 <= msg_in_19; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_20 <= 0; else msg_out_20 <= msg_in_20; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_21 <= 0; else msg_out_21 <= msg_in_21; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_22 <= 0; else msg_out_22 <= msg_in_22; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_23 <= 0; else msg_out_23 <= msg_in_23; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_24 <= 0; else msg_out_24 <= msg_in_24; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_25 <= 0; else msg_out_25 <= msg_in_25; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_26 <= 0; else msg_out_26 <= msg_in_26; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_27 <= 0; else msg_out_27 <= msg_in_27; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_28 <= 0; else msg_out_28 <= msg_in_28; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_29 <= 0; else msg_out_29 <= msg_in_29; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_30 <= 0; else msg_out_30 <= msg_in_30; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_31 <= 0; else msg_out_31 <= msg_in_31; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_32 <= 0; else msg_out_32 <= msg_in_32; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_33 <= 0; else msg_out_33 <= msg_in_33; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_34 <= 0; else msg_out_34 <= msg_in_34; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_35 <= 0; else msg_out_35 <= msg_in_35; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_36 <= 0; else msg_out_36 <= msg_in_36; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_37 <= 0; else msg_out_37 <= msg_in_37; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_38 <= 0; else msg_out_38 <= msg_in_38; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_39 <= 0; else msg_out_39 <= msg_in_39; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_40 <= 0; else msg_out_40 <= msg_in_40; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_41 <= 0; else msg_out_41 <= msg_in_41; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_42 <= 0; else msg_out_42 <= msg_in_42; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_43 <= 0; else msg_out_43 <= msg_in_43; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_44 <= 0; else msg_out_44 <= msg_in_44; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_45 <= 0; else msg_out_45 <= msg_in_45; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_46 <= 0; else msg_out_46 <= msg_in_46; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_47 <= 0; else msg_out_47 <= msg_in_47; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_48 <= 0; else msg_out_48 <= msg_in_48; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_49 <= 0; else msg_out_49 <= msg_in_49; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_50 <= 0; else msg_out_50 <= msg_in_50; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_51 <= 0; else msg_out_51 <= msg_in_51; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_52 <= 0; else msg_out_52 <= msg_in_52; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_53 <= 0; else msg_out_53 <= msg_in_53; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_54 <= 0; else msg_out_54 <= msg_in_54; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_55 <= 0; else msg_out_55 <= msg_in_55; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_56 <= 0; else msg_out_56 <= msg_in_56; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_57 <= 0; else msg_out_57 <= msg_in_57; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_58 <= 0; else msg_out_58 <= msg_in_58; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_59 <= 0; else msg_out_59 <= msg_in_59; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_60 <= 0; else msg_out_60 <= msg_in_60; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_61 <= 0; else msg_out_61 <= msg_in_61; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_62 <= 0; else msg_out_62 <= msg_in_62; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_63 <= 0; else msg_out_63 <= msg_in_63; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_64 <= 0; else msg_out_64 <= msg_in_64; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_65 <= 0; else msg_out_65 <= msg_in_65; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_66 <= 0; else msg_out_66 <= msg_in_66; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_67 <= 0; else msg_out_67 <= msg_in_67; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_68 <= 0; else msg_out_68 <= msg_in_68; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_69 <= 0; else msg_out_69 <= msg_in_69; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_70 <= 0; else msg_out_70 <= msg_in_70; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_71 <= 0; else msg_out_71 <= msg_in_71; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_72 <= 0; else msg_out_72 <= msg_in_72; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_73 <= 0; else msg_out_73 <= msg_in_73; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_74 <= 0; else msg_out_74 <= msg_in_74; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_75 <= 0; else msg_out_75 <= msg_in_75; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_76 <= 0; else msg_out_76 <= msg_in_76; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_77 <= 0; else msg_out_77 <= msg_in_77; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_78 <= 0; else msg_out_78 <= msg_in_78; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_79 <= 0; else msg_out_79 <= msg_in_79; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_80 <= 0; else msg_out_80 <= msg_in_80; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_81 <= 0; else msg_out_81 <= msg_in_81; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_82 <= 0; else msg_out_82 <= msg_in_82; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_83 <= 0; else msg_out_83 <= msg_in_83; end
always @(posedge sys_clk) begin if(rstn == 1'b0) msg_out_84 <= 0; else msg_out_84 <= msg_in_84; end
endmodule
`endif