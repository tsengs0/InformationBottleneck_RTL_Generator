`include "define.vh"

`ifdef SCHED_4_6
module parital_mem_subsystem_top_submatrix_1_3_5_7_9 #(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 255,
	parameter LAYER_NUM = 3,
	parameter CH_DATA_WIDTH = CHECK_PARALLELISM*QUAN_SIZE,
	// Parameters of extrinsic RAMs
	parameter RAM_PORTA_RANGE = 28, // 28 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port A,
	parameter RAM_PORTB_RANGE = 28, // 28 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port b, 
	parameter MEM_DEVICE_NUM = 28,
	parameter DEPTH = 1024,
	parameter DATA_WIDTH = 36,
	parameter FRAG_DATA_WIDTH = 12,
	parameter ADDR_WIDTH = $clog2(DEPTH)
) (
	output wire [CHECK_PARALLELISM-1:0] vnu_pa_msg_bit0,
	output wire [CH_DATA_WIDTH-1:0] pa_to_ch_ram,
	// The memory Dout port to variable nodes as instrinsic messages
	output wire [QUAN_SIZE-1:0] mem_to_vnu_0,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_1,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_2,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_3,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_4,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_5,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_6,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_7,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_8,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_9,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_10,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_11,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_12,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_13,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_14,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_15,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_16,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_17,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_18,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_19,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_20,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_21,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_22,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_23,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_24,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_25,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_26,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_27,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_28,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_29,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_30,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_31,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_32,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_33,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_34,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_35,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_36,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_37,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_38,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_39,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_40,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_41,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_42,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_43,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_44,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_45,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_46,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_47,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_48,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_49,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_50,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_51,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_52,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_53,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_54,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_55,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_56,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_57,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_58,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_59,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_60,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_61,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_62,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_63,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_64,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_65,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_66,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_67,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_68,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_69,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_70,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_71,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_72,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_73,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_74,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_75,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_76,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_77,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_78,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_79,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_80,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_81,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_82,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_83,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_84,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_85,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_86,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_87,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_88,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_89,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_90,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_91,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_92,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_93,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_94,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_95,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_96,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_97,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_98,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_99,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_100,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_101,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_102,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_103,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_104,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_105,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_106,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_107,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_108,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_109,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_110,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_111,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_112,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_113,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_114,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_115,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_116,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_117,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_118,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_119,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_120,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_121,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_122,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_123,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_124,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_125,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_126,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_127,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_128,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_129,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_130,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_131,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_132,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_133,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_134,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_135,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_136,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_137,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_138,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_139,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_140,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_141,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_142,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_143,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_144,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_145,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_146,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_147,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_148,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_149,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_150,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_151,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_152,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_153,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_154,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_155,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_156,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_157,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_158,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_159,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_160,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_161,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_162,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_163,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_164,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_165,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_166,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_167,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_168,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_169,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_170,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_171,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_172,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_173,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_174,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_175,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_176,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_177,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_178,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_179,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_180,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_181,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_182,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_183,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_184,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_185,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_186,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_187,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_188,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_189,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_190,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_191,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_192,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_193,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_194,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_195,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_196,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_197,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_198,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_199,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_200,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_201,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_202,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_203,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_204,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_205,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_206,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_207,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_208,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_209,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_210,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_211,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_212,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_213,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_214,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_215,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_216,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_217,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_218,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_219,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_220,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_221,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_222,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_223,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_224,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_225,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_226,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_227,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_228,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_229,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_230,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_231,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_232,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_233,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_234,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_235,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_236,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_237,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_238,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_239,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_240,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_241,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_242,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_243,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_244,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_245,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_246,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_247,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_248,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_249,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_250,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_251,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_252,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_253,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_254,
	// The memory Dout port to check nodes as instrinsic messages
	output wire [QUAN_SIZE-1:0] mem_to_cnu_0,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_1,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_2,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_3,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_4,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_5,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_6,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_7,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_8,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_9,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_10,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_11,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_12,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_13,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_14,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_15,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_16,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_17,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_18,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_19,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_20,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_21,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_22,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_23,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_24,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_25,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_26,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_27,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_28,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_29,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_30,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_31,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_32,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_33,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_34,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_35,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_36,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_37,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_38,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_39,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_40,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_41,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_42,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_43,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_44,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_45,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_46,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_47,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_48,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_49,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_50,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_51,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_52,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_53,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_54,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_55,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_56,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_57,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_58,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_59,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_60,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_61,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_62,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_63,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_64,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_65,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_66,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_67,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_68,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_69,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_70,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_71,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_72,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_73,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_74,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_75,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_76,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_77,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_78,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_79,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_80,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_81,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_82,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_83,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_84,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_85,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_86,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_87,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_88,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_89,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_90,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_91,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_92,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_93,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_94,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_95,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_96,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_97,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_98,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_99,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_100,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_101,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_102,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_103,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_104,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_105,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_106,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_107,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_108,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_109,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_110,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_111,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_112,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_113,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_114,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_115,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_116,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_117,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_118,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_119,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_120,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_121,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_122,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_123,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_124,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_125,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_126,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_127,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_128,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_129,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_130,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_131,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_132,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_133,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_134,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_135,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_136,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_137,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_138,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_139,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_140,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_141,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_142,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_143,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_144,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_145,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_146,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_147,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_148,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_149,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_150,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_151,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_152,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_153,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_154,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_155,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_156,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_157,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_158,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_159,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_160,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_161,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_162,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_163,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_164,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_165,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_166,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_167,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_168,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_169,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_170,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_171,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_172,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_173,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_174,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_175,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_176,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_177,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_178,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_179,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_180,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_181,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_182,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_183,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_184,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_185,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_186,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_187,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_188,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_189,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_190,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_191,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_192,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_193,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_194,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_195,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_196,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_197,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_198,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_199,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_200,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_201,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_202,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_203,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_204,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_205,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_206,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_207,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_208,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_209,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_210,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_211,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_212,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_213,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_214,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_215,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_216,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_217,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_218,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_219,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_220,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_221,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_222,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_223,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_224,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_225,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_226,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_227,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_228,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_229,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_230,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_231,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_232,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_233,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_234,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_235,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_236,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_237,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_238,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_239,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_240,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_241,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_242,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_243,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_244,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_245,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_246,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_247,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_248,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_249,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_250,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_251,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_252,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_253,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_254,
	// The varible extrinsic message written back onto memory through BS and PA
	input wire [QUAN_SIZE-1:0] vnu_to_mem_0,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_1,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_2,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_3,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_4,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_5,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_6,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_7,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_8,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_9,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_10,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_11,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_12,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_13,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_14,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_15,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_16,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_17,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_18,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_19,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_20,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_21,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_22,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_23,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_24,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_25,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_26,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_27,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_28,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_29,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_30,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_31,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_32,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_33,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_34,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_35,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_36,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_37,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_38,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_39,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_40,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_41,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_42,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_43,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_44,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_45,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_46,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_47,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_48,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_49,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_50,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_51,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_52,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_53,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_54,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_55,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_56,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_57,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_58,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_59,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_60,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_61,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_62,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_63,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_64,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_65,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_66,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_67,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_68,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_69,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_70,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_71,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_72,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_73,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_74,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_75,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_76,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_77,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_78,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_79,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_80,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_81,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_82,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_83,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_84,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_85,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_86,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_87,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_88,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_89,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_90,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_91,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_92,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_93,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_94,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_95,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_96,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_97,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_98,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_99,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_100,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_101,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_102,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_103,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_104,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_105,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_106,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_107,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_108,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_109,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_110,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_111,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_112,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_113,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_114,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_115,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_116,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_117,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_118,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_119,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_120,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_121,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_122,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_123,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_124,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_125,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_126,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_127,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_128,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_129,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_130,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_131,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_132,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_133,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_134,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_135,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_136,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_137,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_138,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_139,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_140,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_141,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_142,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_143,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_144,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_145,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_146,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_147,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_148,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_149,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_150,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_151,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_152,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_153,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_154,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_155,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_156,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_157,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_158,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_159,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_160,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_161,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_162,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_163,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_164,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_165,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_166,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_167,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_168,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_169,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_170,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_171,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_172,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_173,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_174,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_175,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_176,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_177,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_178,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_179,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_180,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_181,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_182,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_183,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_184,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_185,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_186,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_187,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_188,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_189,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_190,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_191,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_192,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_193,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_194,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_195,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_196,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_197,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_198,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_199,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_200,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_201,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_202,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_203,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_204,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_205,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_206,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_207,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_208,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_209,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_210,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_211,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_212,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_213,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_214,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_215,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_216,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_217,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_218,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_219,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_220,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_221,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_222,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_223,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_224,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_225,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_226,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_227,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_228,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_229,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_230,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_231,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_232,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_233,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_234,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_235,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_236,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_237,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_238,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_239,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_240,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_241,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_242,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_243,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_244,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_245,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_246,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_247,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_248,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_249,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_250,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_251,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_252,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_253,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_254,
	// The check extrinsic message written back onto memory through BS and PA
	input wire [QUAN_SIZE-1:0] cnu_to_mem_0,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_1,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_2,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_3,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_4,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_5,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_6,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_7,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_8,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_9,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_10,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_11,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_12,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_13,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_14,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_15,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_16,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_17,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_18,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_19,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_20,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_21,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_22,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_23,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_24,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_25,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_26,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_27,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_28,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_29,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_30,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_31,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_32,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_33,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_34,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_35,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_36,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_37,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_38,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_39,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_40,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_41,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_42,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_43,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_44,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_45,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_46,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_47,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_48,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_49,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_50,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_51,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_52,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_53,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_54,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_55,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_56,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_57,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_58,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_59,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_60,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_61,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_62,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_63,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_64,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_65,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_66,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_67,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_68,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_69,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_70,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_71,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_72,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_73,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_74,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_75,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_76,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_77,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_78,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_79,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_80,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_81,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_82,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_83,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_84,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_85,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_86,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_87,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_88,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_89,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_90,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_91,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_92,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_93,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_94,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_95,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_96,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_97,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_98,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_99,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_100,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_101,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_102,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_103,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_104,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_105,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_106,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_107,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_108,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_109,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_110,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_111,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_112,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_113,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_114,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_115,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_116,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_117,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_118,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_119,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_120,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_121,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_122,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_123,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_124,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_125,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_126,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_127,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_128,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_129,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_130,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_131,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_132,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_133,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_134,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_135,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_136,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_137,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_138,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_139,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_140,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_141,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_142,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_143,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_144,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_145,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_146,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_147,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_148,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_149,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_150,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_151,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_152,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_153,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_154,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_155,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_156,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_157,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_158,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_159,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_160,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_161,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_162,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_163,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_164,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_165,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_166,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_167,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_168,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_169,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_170,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_171,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_172,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_173,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_174,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_175,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_176,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_177,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_178,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_179,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_180,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_181,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_182,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_183,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_184,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_185,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_186,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_187,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_188,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_189,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_190,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_191,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_192,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_193,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_194,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_195,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_196,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_197,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_198,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_199,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_200,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_201,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_202,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_203,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_204,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_205,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_206,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_207,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_208,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_209,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_210,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_211,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_212,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_213,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_214,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_215,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_216,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_217,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_218,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_219,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_220,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_221,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_222,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_223,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_224,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_225,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_226,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_227,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_228,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_229,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_230,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_231,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_232,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_233,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_234,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_235,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_236,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_237,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_238,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_239,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_240,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_241,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_242,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_243,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_244,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_245,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_246,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_247,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_248,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_249,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_250,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_251,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_252,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_253,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_254,

	input wire [ADDR_WIDTH-1:0] cnu_sync_addr,
	input wire [ADDR_WIDTH-1:0] vnu_sync_addr,
	input wire [LAYER_NUM-1:0] cnu_layer_status,
	input wire [LAYER_NUM-1:0] vnu_layer_status,
	input wire [`ROW_SPLIT_FACTOR-1:0] cnu_sub_row_status,
	input wire [`ROW_SPLIT_FACTOR-1:0] vnu_sub_row_status,
	input wire [1:0] last_row_chunk, // [0]: check; [1]: variable
	input wire [1:0] we, // [0]: check; [1]: variable
	input wire sys_clk,
	input wire rstn
);
/*-------------------------------------------------------*/
// Page alignment of Check nodes
wire [QUAN_SIZE-1:0] cnu_pa_msg [CHECK_PARALLELISM-1:0];
ram_pageAlign_interface_partial_col_1_3_5_7_9 #(
	.QUAN_SIZE(QUAN_SIZE),
	.CHECK_PARALLELISM(CHECK_PARALLELISM),
	.LAYER_NUM(LAYER_NUM)
) cnu_ram_pageAlign_interface_submatrix_1_3_5_7_9 (
	.msg_out_0			(cnu_pa_msg[0]),
	.msg_out_1			(cnu_pa_msg[1]),
	.msg_out_2			(cnu_pa_msg[2]),
	.msg_out_3			(cnu_pa_msg[3]),
	.msg_out_4			(cnu_pa_msg[4]),
	.msg_out_5			(cnu_pa_msg[5]),
	.msg_out_6			(cnu_pa_msg[6]),
	.msg_out_7			(cnu_pa_msg[7]),
	.msg_out_8			(cnu_pa_msg[8]),
	.msg_out_9			(cnu_pa_msg[9]),
	.msg_out_10			(cnu_pa_msg[10]),
	.msg_out_11			(cnu_pa_msg[11]),
	.msg_out_12			(cnu_pa_msg[12]),
	.msg_out_13			(cnu_pa_msg[13]),
	.msg_out_14			(cnu_pa_msg[14]),
	.msg_out_15			(cnu_pa_msg[15]),
	.msg_out_16			(cnu_pa_msg[16]),
	.msg_out_17			(cnu_pa_msg[17]),
	.msg_out_18			(cnu_pa_msg[18]),
	.msg_out_19			(cnu_pa_msg[19]),
	.msg_out_20			(cnu_pa_msg[20]),
	.msg_out_21			(cnu_pa_msg[21]),
	.msg_out_22			(cnu_pa_msg[22]),
	.msg_out_23			(cnu_pa_msg[23]),
	.msg_out_24			(cnu_pa_msg[24]),
	.msg_out_25			(cnu_pa_msg[25]),
	.msg_out_26			(cnu_pa_msg[26]),
	.msg_out_27			(cnu_pa_msg[27]),
	.msg_out_28			(cnu_pa_msg[28]),
	.msg_out_29			(cnu_pa_msg[29]),
	.msg_out_30			(cnu_pa_msg[30]),
	.msg_out_31			(cnu_pa_msg[31]),
	.msg_out_32			(cnu_pa_msg[32]),
	.msg_out_33			(cnu_pa_msg[33]),
	.msg_out_34			(cnu_pa_msg[34]),
	.msg_out_35			(cnu_pa_msg[35]),
	.msg_out_36			(cnu_pa_msg[36]),
	.msg_out_37			(cnu_pa_msg[37]),
	.msg_out_38			(cnu_pa_msg[38]),
	.msg_out_39			(cnu_pa_msg[39]),
	.msg_out_40			(cnu_pa_msg[40]),
	.msg_out_41			(cnu_pa_msg[41]),
	.msg_out_42			(cnu_pa_msg[42]),
	.msg_out_43			(cnu_pa_msg[43]),
	.msg_out_44			(cnu_pa_msg[44]),
	.msg_out_45			(cnu_pa_msg[45]),
	.msg_out_46			(cnu_pa_msg[46]),
	.msg_out_47			(cnu_pa_msg[47]),
	.msg_out_48			(cnu_pa_msg[48]),
	.msg_out_49			(cnu_pa_msg[49]),
	.msg_out_50			(cnu_pa_msg[50]),
	.msg_out_51			(cnu_pa_msg[51]),
	.msg_out_52			(cnu_pa_msg[52]),
	.msg_out_53			(cnu_pa_msg[53]),
	.msg_out_54			(cnu_pa_msg[54]),
	.msg_out_55			(cnu_pa_msg[55]),
	.msg_out_56			(cnu_pa_msg[56]),
	.msg_out_57			(cnu_pa_msg[57]),
	.msg_out_58			(cnu_pa_msg[58]),
	.msg_out_59			(cnu_pa_msg[59]),
	.msg_out_60			(cnu_pa_msg[60]),
	.msg_out_61			(cnu_pa_msg[61]),
	.msg_out_62			(cnu_pa_msg[62]),
	.msg_out_63			(cnu_pa_msg[63]),
	.msg_out_64			(cnu_pa_msg[64]),
	.msg_out_65			(cnu_pa_msg[65]),
	.msg_out_66			(cnu_pa_msg[66]),
	.msg_out_67			(cnu_pa_msg[67]),
	.msg_out_68			(cnu_pa_msg[68]),
	.msg_out_69			(cnu_pa_msg[69]),
	.msg_out_70			(cnu_pa_msg[70]),
	.msg_out_71			(cnu_pa_msg[71]),
	.msg_out_72			(cnu_pa_msg[72]),
	.msg_out_73			(cnu_pa_msg[73]),
	.msg_out_74			(cnu_pa_msg[74]),
	.msg_out_75			(cnu_pa_msg[75]),
	.msg_out_76			(cnu_pa_msg[76]),
	.msg_out_77			(cnu_pa_msg[77]),
	.msg_out_78			(cnu_pa_msg[78]),
	.msg_out_79			(cnu_pa_msg[79]),
	.msg_out_80			(cnu_pa_msg[80]),
	.msg_out_81			(cnu_pa_msg[81]),
	.msg_out_82			(cnu_pa_msg[82]),
	.msg_out_83			(cnu_pa_msg[83]),
	.msg_out_84			(cnu_pa_msg[84]),
	.msg_out_85			(cnu_pa_msg[85]),
	.msg_out_86			(cnu_pa_msg[86]),
	.msg_out_87			(cnu_pa_msg[87]),
	.msg_out_88			(cnu_pa_msg[88]),
	.msg_out_89			(cnu_pa_msg[89]),
	.msg_out_90			(cnu_pa_msg[90]),
	.msg_out_91			(cnu_pa_msg[91]),
	.msg_out_92			(cnu_pa_msg[92]),
	.msg_out_93			(cnu_pa_msg[93]),
	.msg_out_94			(cnu_pa_msg[94]),
	.msg_out_95			(cnu_pa_msg[95]),
	.msg_out_96			(cnu_pa_msg[96]),
	.msg_out_97			(cnu_pa_msg[97]),
	.msg_out_98			(cnu_pa_msg[98]),
	.msg_out_99			(cnu_pa_msg[99]),
	.msg_out_100			(cnu_pa_msg[100]),
	.msg_out_101			(cnu_pa_msg[101]),
	.msg_out_102			(cnu_pa_msg[102]),
	.msg_out_103			(cnu_pa_msg[103]),
	.msg_out_104			(cnu_pa_msg[104]),
	.msg_out_105			(cnu_pa_msg[105]),
	.msg_out_106			(cnu_pa_msg[106]),
	.msg_out_107			(cnu_pa_msg[107]),
	.msg_out_108			(cnu_pa_msg[108]),
	.msg_out_109			(cnu_pa_msg[109]),
	.msg_out_110			(cnu_pa_msg[110]),
	.msg_out_111			(cnu_pa_msg[111]),
	.msg_out_112			(cnu_pa_msg[112]),
	.msg_out_113			(cnu_pa_msg[113]),
	.msg_out_114			(cnu_pa_msg[114]),
	.msg_out_115			(cnu_pa_msg[115]),
	.msg_out_116			(cnu_pa_msg[116]),
	.msg_out_117			(cnu_pa_msg[117]),
	.msg_out_118			(cnu_pa_msg[118]),
	.msg_out_119			(cnu_pa_msg[119]),
	.msg_out_120			(cnu_pa_msg[120]),
	.msg_out_121			(cnu_pa_msg[121]),
	.msg_out_122			(cnu_pa_msg[122]),
	.msg_out_123			(cnu_pa_msg[123]),
	.msg_out_124			(cnu_pa_msg[124]),
	.msg_out_125			(cnu_pa_msg[125]),
	.msg_out_126			(cnu_pa_msg[126]),
	.msg_out_127			(cnu_pa_msg[127]),
	.msg_out_128			(cnu_pa_msg[128]),
	.msg_out_129			(cnu_pa_msg[129]),
	.msg_out_130			(cnu_pa_msg[130]),
	.msg_out_131			(cnu_pa_msg[131]),
	.msg_out_132			(cnu_pa_msg[132]),
	.msg_out_133			(cnu_pa_msg[133]),
	.msg_out_134			(cnu_pa_msg[134]),
	.msg_out_135			(cnu_pa_msg[135]),
	.msg_out_136			(cnu_pa_msg[136]),
	.msg_out_137			(cnu_pa_msg[137]),
	.msg_out_138			(cnu_pa_msg[138]),
	.msg_out_139			(cnu_pa_msg[139]),
	.msg_out_140			(cnu_pa_msg[140]),
	.msg_out_141			(cnu_pa_msg[141]),
	.msg_out_142			(cnu_pa_msg[142]),
	.msg_out_143			(cnu_pa_msg[143]),
	.msg_out_144			(cnu_pa_msg[144]),
	.msg_out_145			(cnu_pa_msg[145]),
	.msg_out_146			(cnu_pa_msg[146]),
	.msg_out_147			(cnu_pa_msg[147]),
	.msg_out_148			(cnu_pa_msg[148]),
	.msg_out_149			(cnu_pa_msg[149]),
	.msg_out_150			(cnu_pa_msg[150]),
	.msg_out_151			(cnu_pa_msg[151]),
	.msg_out_152			(cnu_pa_msg[152]),
	.msg_out_153			(cnu_pa_msg[153]),
	.msg_out_154			(cnu_pa_msg[154]),
	.msg_out_155			(cnu_pa_msg[155]),
	.msg_out_156			(cnu_pa_msg[156]),
	.msg_out_157			(cnu_pa_msg[157]),
	.msg_out_158			(cnu_pa_msg[158]),
	.msg_out_159			(cnu_pa_msg[159]),
	.msg_out_160			(cnu_pa_msg[160]),
	.msg_out_161			(cnu_pa_msg[161]),
	.msg_out_162			(cnu_pa_msg[162]),
	.msg_out_163			(cnu_pa_msg[163]),
	.msg_out_164			(cnu_pa_msg[164]),
	.msg_out_165			(cnu_pa_msg[165]),
	.msg_out_166			(cnu_pa_msg[166]),
	.msg_out_167			(cnu_pa_msg[167]),
	.msg_out_168			(cnu_pa_msg[168]),
	.msg_out_169			(cnu_pa_msg[169]),
	.msg_out_170			(cnu_pa_msg[170]),
	.msg_out_171			(cnu_pa_msg[171]),
	.msg_out_172			(cnu_pa_msg[172]),
	.msg_out_173			(cnu_pa_msg[173]),
	.msg_out_174			(cnu_pa_msg[174]),
	.msg_out_175			(cnu_pa_msg[175]),
	.msg_out_176			(cnu_pa_msg[176]),
	.msg_out_177			(cnu_pa_msg[177]),
	.msg_out_178			(cnu_pa_msg[178]),
	.msg_out_179			(cnu_pa_msg[179]),
	.msg_out_180			(cnu_pa_msg[180]),
	.msg_out_181			(cnu_pa_msg[181]),
	.msg_out_182			(cnu_pa_msg[182]),
	.msg_out_183			(cnu_pa_msg[183]),
	.msg_out_184			(cnu_pa_msg[184]),
	.msg_out_185			(cnu_pa_msg[185]),
	.msg_out_186			(cnu_pa_msg[186]),
	.msg_out_187			(cnu_pa_msg[187]),
	.msg_out_188			(cnu_pa_msg[188]),
	.msg_out_189			(cnu_pa_msg[189]),
	.msg_out_190			(cnu_pa_msg[190]),
	.msg_out_191			(cnu_pa_msg[191]),
	.msg_out_192			(cnu_pa_msg[192]),
	.msg_out_193			(cnu_pa_msg[193]),
	.msg_out_194			(cnu_pa_msg[194]),
	.msg_out_195			(cnu_pa_msg[195]),
	.msg_out_196			(cnu_pa_msg[196]),
	.msg_out_197			(cnu_pa_msg[197]),
	.msg_out_198			(cnu_pa_msg[198]),
	.msg_out_199			(cnu_pa_msg[199]),
	.msg_out_200			(cnu_pa_msg[200]),
	.msg_out_201			(cnu_pa_msg[201]),
	.msg_out_202			(cnu_pa_msg[202]),
	.msg_out_203			(cnu_pa_msg[203]),
	.msg_out_204			(cnu_pa_msg[204]),
	.msg_out_205			(cnu_pa_msg[205]),
	.msg_out_206			(cnu_pa_msg[206]),
	.msg_out_207			(cnu_pa_msg[207]),
	.msg_out_208			(cnu_pa_msg[208]),
	.msg_out_209			(cnu_pa_msg[209]),
	.msg_out_210			(cnu_pa_msg[210]),
	.msg_out_211			(cnu_pa_msg[211]),
	.msg_out_212			(cnu_pa_msg[212]),
	.msg_out_213			(cnu_pa_msg[213]),
	.msg_out_214			(cnu_pa_msg[214]),
	.msg_out_215			(cnu_pa_msg[215]),
	.msg_out_216			(cnu_pa_msg[216]),
	.msg_out_217			(cnu_pa_msg[217]),
	.msg_out_218			(cnu_pa_msg[218]),
	.msg_out_219			(cnu_pa_msg[219]),
	.msg_out_220			(cnu_pa_msg[220]),
	.msg_out_221			(cnu_pa_msg[221]),
	.msg_out_222			(cnu_pa_msg[222]),
	.msg_out_223			(cnu_pa_msg[223]),
	.msg_out_224			(cnu_pa_msg[224]),
	.msg_out_225			(cnu_pa_msg[225]),
	.msg_out_226			(cnu_pa_msg[226]),
	.msg_out_227			(cnu_pa_msg[227]),
	.msg_out_228			(cnu_pa_msg[228]),
	.msg_out_229			(cnu_pa_msg[229]),
	.msg_out_230			(cnu_pa_msg[230]),
	.msg_out_231			(cnu_pa_msg[231]),
	.msg_out_232			(cnu_pa_msg[232]),
	.msg_out_233			(cnu_pa_msg[233]),
	.msg_out_234			(cnu_pa_msg[234]),
	.msg_out_235			(cnu_pa_msg[235]),
	.msg_out_236			(cnu_pa_msg[236]),
	.msg_out_237			(cnu_pa_msg[237]),
	.msg_out_238			(cnu_pa_msg[238]),
	.msg_out_239			(cnu_pa_msg[239]),
	.msg_out_240			(cnu_pa_msg[240]),
	.msg_out_241			(cnu_pa_msg[241]),
	.msg_out_242			(cnu_pa_msg[242]),
	.msg_out_243			(cnu_pa_msg[243]),
	.msg_out_244			(cnu_pa_msg[244]),
	.msg_out_245			(cnu_pa_msg[245]),
	.msg_out_246			(cnu_pa_msg[246]),
	.msg_out_247			(cnu_pa_msg[247]),
	.msg_out_248			(cnu_pa_msg[248]),
	.msg_out_249			(cnu_pa_msg[249]),
	.msg_out_250			(cnu_pa_msg[250]),
	.msg_out_251			(cnu_pa_msg[251]),
	.msg_out_252			(cnu_pa_msg[252]),
	.msg_out_253			(cnu_pa_msg[253]),
	.msg_out_254			(cnu_pa_msg[254]),
	.msg_in_0			(cnu_to_mem_0),
	.msg_in_1			(cnu_to_mem_1),
	.msg_in_2			(cnu_to_mem_2),
	.msg_in_3			(cnu_to_mem_3),
	.msg_in_4			(cnu_to_mem_4),
	.msg_in_5			(cnu_to_mem_5),
	.msg_in_6			(cnu_to_mem_6),
	.msg_in_7			(cnu_to_mem_7),
	.msg_in_8			(cnu_to_mem_8),
	.msg_in_9			(cnu_to_mem_9),
	.msg_in_10			(cnu_to_mem_10),
	.msg_in_11			(cnu_to_mem_11),
	.msg_in_12			(cnu_to_mem_12),
	.msg_in_13			(cnu_to_mem_13),
	.msg_in_14			(cnu_to_mem_14),
	.msg_in_15			(cnu_to_mem_15),
	.msg_in_16			(cnu_to_mem_16),
	.msg_in_17			(cnu_to_mem_17),
	.msg_in_18			(cnu_to_mem_18),
	.msg_in_19			(cnu_to_mem_19),
	.msg_in_20			(cnu_to_mem_20),
	.msg_in_21			(cnu_to_mem_21),
	.msg_in_22			(cnu_to_mem_22),
	.msg_in_23			(cnu_to_mem_23),
	.msg_in_24			(cnu_to_mem_24),
	.msg_in_25			(cnu_to_mem_25),
	.msg_in_26			(cnu_to_mem_26),
	.msg_in_27			(cnu_to_mem_27),
	.msg_in_28			(cnu_to_mem_28),
	.msg_in_29			(cnu_to_mem_29),
	.msg_in_30			(cnu_to_mem_30),
	.msg_in_31			(cnu_to_mem_31),
	.msg_in_32			(cnu_to_mem_32),
	.msg_in_33			(cnu_to_mem_33),
	.msg_in_34			(cnu_to_mem_34),
	.msg_in_35			(cnu_to_mem_35),
	.msg_in_36			(cnu_to_mem_36),
	.msg_in_37			(cnu_to_mem_37),
	.msg_in_38			(cnu_to_mem_38),
	.msg_in_39			(cnu_to_mem_39),
	.msg_in_40			(cnu_to_mem_40),
	.msg_in_41			(cnu_to_mem_41),
	.msg_in_42			(cnu_to_mem_42),
	.msg_in_43			(cnu_to_mem_43),
	.msg_in_44			(cnu_to_mem_44),
	.msg_in_45			(cnu_to_mem_45),
	.msg_in_46			(cnu_to_mem_46),
	.msg_in_47			(cnu_to_mem_47),
	.msg_in_48			(cnu_to_mem_48),
	.msg_in_49			(cnu_to_mem_49),
	.msg_in_50			(cnu_to_mem_50),
	.msg_in_51			(cnu_to_mem_51),
	.msg_in_52			(cnu_to_mem_52),
	.msg_in_53			(cnu_to_mem_53),
	.msg_in_54			(cnu_to_mem_54),
	.msg_in_55			(cnu_to_mem_55),
	.msg_in_56			(cnu_to_mem_56),
	.msg_in_57			(cnu_to_mem_57),
	.msg_in_58			(cnu_to_mem_58),
	.msg_in_59			(cnu_to_mem_59),
	.msg_in_60			(cnu_to_mem_60),
	.msg_in_61			(cnu_to_mem_61),
	.msg_in_62			(cnu_to_mem_62),
	.msg_in_63			(cnu_to_mem_63),
	.msg_in_64			(cnu_to_mem_64),
	.msg_in_65			(cnu_to_mem_65),
	.msg_in_66			(cnu_to_mem_66),
	.msg_in_67			(cnu_to_mem_67),
	.msg_in_68			(cnu_to_mem_68),
	.msg_in_69			(cnu_to_mem_69),
	.msg_in_70			(cnu_to_mem_70),
	.msg_in_71			(cnu_to_mem_71),
	.msg_in_72			(cnu_to_mem_72),
	.msg_in_73			(cnu_to_mem_73),
	.msg_in_74			(cnu_to_mem_74),
	.msg_in_75			(cnu_to_mem_75),
	.msg_in_76			(cnu_to_mem_76),
	.msg_in_77			(cnu_to_mem_77),
	.msg_in_78			(cnu_to_mem_78),
	.msg_in_79			(cnu_to_mem_79),
	.msg_in_80			(cnu_to_mem_80),
	.msg_in_81			(cnu_to_mem_81),
	.msg_in_82			(cnu_to_mem_82),
	.msg_in_83			(cnu_to_mem_83),
	.msg_in_84			(cnu_to_mem_84),
	.msg_in_85			(cnu_to_mem_85),
	.msg_in_86			(cnu_to_mem_86),
	.msg_in_87			(cnu_to_mem_87),
	.msg_in_88			(cnu_to_mem_88),
	.msg_in_89			(cnu_to_mem_89),
	.msg_in_90			(cnu_to_mem_90),
	.msg_in_91			(cnu_to_mem_91),
	.msg_in_92			(cnu_to_mem_92),
	.msg_in_93			(cnu_to_mem_93),
	.msg_in_94			(cnu_to_mem_94),
	.msg_in_95			(cnu_to_mem_95),
	.msg_in_96			(cnu_to_mem_96),
	.msg_in_97			(cnu_to_mem_97),
	.msg_in_98			(cnu_to_mem_98),
	.msg_in_99			(cnu_to_mem_99),
	.msg_in_100			(cnu_to_mem_100),
	.msg_in_101			(cnu_to_mem_101),
	.msg_in_102			(cnu_to_mem_102),
	.msg_in_103			(cnu_to_mem_103),
	.msg_in_104			(cnu_to_mem_104),
	.msg_in_105			(cnu_to_mem_105),
	.msg_in_106			(cnu_to_mem_106),
	.msg_in_107			(cnu_to_mem_107),
	.msg_in_108			(cnu_to_mem_108),
	.msg_in_109			(cnu_to_mem_109),
	.msg_in_110			(cnu_to_mem_110),
	.msg_in_111			(cnu_to_mem_111),
	.msg_in_112			(cnu_to_mem_112),
	.msg_in_113			(cnu_to_mem_113),
	.msg_in_114			(cnu_to_mem_114),
	.msg_in_115			(cnu_to_mem_115),
	.msg_in_116			(cnu_to_mem_116),
	.msg_in_117			(cnu_to_mem_117),
	.msg_in_118			(cnu_to_mem_118),
	.msg_in_119			(cnu_to_mem_119),
	.msg_in_120			(cnu_to_mem_120),
	.msg_in_121			(cnu_to_mem_121),
	.msg_in_122			(cnu_to_mem_122),
	.msg_in_123			(cnu_to_mem_123),
	.msg_in_124			(cnu_to_mem_124),
	.msg_in_125			(cnu_to_mem_125),
	.msg_in_126			(cnu_to_mem_126),
	.msg_in_127			(cnu_to_mem_127),
	.msg_in_128			(cnu_to_mem_128),
	.msg_in_129			(cnu_to_mem_129),
	.msg_in_130			(cnu_to_mem_130),
	.msg_in_131			(cnu_to_mem_131),
	.msg_in_132			(cnu_to_mem_132),
	.msg_in_133			(cnu_to_mem_133),
	.msg_in_134			(cnu_to_mem_134),
	.msg_in_135			(cnu_to_mem_135),
	.msg_in_136			(cnu_to_mem_136),
	.msg_in_137			(cnu_to_mem_137),
	.msg_in_138			(cnu_to_mem_138),
	.msg_in_139			(cnu_to_mem_139),
	.msg_in_140			(cnu_to_mem_140),
	.msg_in_141			(cnu_to_mem_141),
	.msg_in_142			(cnu_to_mem_142),
	.msg_in_143			(cnu_to_mem_143),
	.msg_in_144			(cnu_to_mem_144),
	.msg_in_145			(cnu_to_mem_145),
	.msg_in_146			(cnu_to_mem_146),
	.msg_in_147			(cnu_to_mem_147),
	.msg_in_148			(cnu_to_mem_148),
	.msg_in_149			(cnu_to_mem_149),
	.msg_in_150			(cnu_to_mem_150),
	.msg_in_151			(cnu_to_mem_151),
	.msg_in_152			(cnu_to_mem_152),
	.msg_in_153			(cnu_to_mem_153),
	.msg_in_154			(cnu_to_mem_154),
	.msg_in_155			(cnu_to_mem_155),
	.msg_in_156			(cnu_to_mem_156),
	.msg_in_157			(cnu_to_mem_157),
	.msg_in_158			(cnu_to_mem_158),
	.msg_in_159			(cnu_to_mem_159),
	.msg_in_160			(cnu_to_mem_160),
	.msg_in_161			(cnu_to_mem_161),
	.msg_in_162			(cnu_to_mem_162),
	.msg_in_163			(cnu_to_mem_163),
	.msg_in_164			(cnu_to_mem_164),
	.msg_in_165			(cnu_to_mem_165),
	.msg_in_166			(cnu_to_mem_166),
	.msg_in_167			(cnu_to_mem_167),
	.msg_in_168			(cnu_to_mem_168),
	.msg_in_169			(cnu_to_mem_169),
	.msg_in_170			(cnu_to_mem_170),
	.msg_in_171			(cnu_to_mem_171),
	.msg_in_172			(cnu_to_mem_172),
	.msg_in_173			(cnu_to_mem_173),
	.msg_in_174			(cnu_to_mem_174),
	.msg_in_175			(cnu_to_mem_175),
	.msg_in_176			(cnu_to_mem_176),
	.msg_in_177			(cnu_to_mem_177),
	.msg_in_178			(cnu_to_mem_178),
	.msg_in_179			(cnu_to_mem_179),
	.msg_in_180			(cnu_to_mem_180),
	.msg_in_181			(cnu_to_mem_181),
	.msg_in_182			(cnu_to_mem_182),
	.msg_in_183			(cnu_to_mem_183),
	.msg_in_184			(cnu_to_mem_184),
	.msg_in_185			(cnu_to_mem_185),
	.msg_in_186			(cnu_to_mem_186),
	.msg_in_187			(cnu_to_mem_187),
	.msg_in_188			(cnu_to_mem_188),
	.msg_in_189			(cnu_to_mem_189),
	.msg_in_190			(cnu_to_mem_190),
	.msg_in_191			(cnu_to_mem_191),
	.msg_in_192			(cnu_to_mem_192),
	.msg_in_193			(cnu_to_mem_193),
	.msg_in_194			(cnu_to_mem_194),
	.msg_in_195			(cnu_to_mem_195),
	.msg_in_196			(cnu_to_mem_196),
	.msg_in_197			(cnu_to_mem_197),
	.msg_in_198			(cnu_to_mem_198),
	.msg_in_199			(cnu_to_mem_199),
	.msg_in_200			(cnu_to_mem_200),
	.msg_in_201			(cnu_to_mem_201),
	.msg_in_202			(cnu_to_mem_202),
	.msg_in_203			(cnu_to_mem_203),
	.msg_in_204			(cnu_to_mem_204),
	.msg_in_205			(cnu_to_mem_205),
	.msg_in_206			(cnu_to_mem_206),
	.msg_in_207			(cnu_to_mem_207),
	.msg_in_208			(cnu_to_mem_208),
	.msg_in_209			(cnu_to_mem_209),
	.msg_in_210			(cnu_to_mem_210),
	.msg_in_211			(cnu_to_mem_211),
	.msg_in_212			(cnu_to_mem_212),
	.msg_in_213			(cnu_to_mem_213),
	.msg_in_214			(cnu_to_mem_214),
	.msg_in_215			(cnu_to_mem_215),
	.msg_in_216			(cnu_to_mem_216),
	.msg_in_217			(cnu_to_mem_217),
	.msg_in_218			(cnu_to_mem_218),
	.msg_in_219			(cnu_to_mem_219),
	.msg_in_220			(cnu_to_mem_220),
	.msg_in_221			(cnu_to_mem_221),
	.msg_in_222			(cnu_to_mem_222),
	.msg_in_223			(cnu_to_mem_223),
	.msg_in_224			(cnu_to_mem_224),
	.msg_in_225			(cnu_to_mem_225),
	.msg_in_226			(cnu_to_mem_226),
	.msg_in_227			(cnu_to_mem_227),
	.msg_in_228			(cnu_to_mem_228),
	.msg_in_229			(cnu_to_mem_229),
	.msg_in_230			(cnu_to_mem_230),
	.msg_in_231			(cnu_to_mem_231),
	.msg_in_232			(cnu_to_mem_232),
	.msg_in_233			(cnu_to_mem_233),
	.msg_in_234			(cnu_to_mem_234),
	.msg_in_235			(cnu_to_mem_235),
	.msg_in_236			(cnu_to_mem_236),
	.msg_in_237			(cnu_to_mem_237),
	.msg_in_238			(cnu_to_mem_238),
	.msg_in_239			(cnu_to_mem_239),
	.msg_in_240			(cnu_to_mem_240),
	.msg_in_241			(cnu_to_mem_241),
	.msg_in_242			(cnu_to_mem_242),
	.msg_in_243			(cnu_to_mem_243),
	.msg_in_244			(cnu_to_mem_244),
	.msg_in_245			(cnu_to_mem_245),
	.msg_in_246			(cnu_to_mem_246),
	.msg_in_247			(cnu_to_mem_247),
	.msg_in_248			(cnu_to_mem_248),
	.msg_in_249			(cnu_to_mem_249),
	.msg_in_250			(cnu_to_mem_250),
	.msg_in_251			(cnu_to_mem_251),
	.msg_in_252			(cnu_to_mem_252),
	.msg_in_253			(cnu_to_mem_253),
	.msg_in_254			(cnu_to_mem_254),
	.layer_status	(cnu_layer_status),
	.first_row_chunk	(last_row_chunk[0]),
	.sub_row_status	(cnu_sub_row_status[`ROW_SPLIT_FACTOR-1:0]),
	.sys_clk	(sys_clk),
	.rstn	(rstn)
);
/*-------------------------------------------------------*/
// Page alignment of Variable nodes
wire [QUAN_SIZE-1:0] vnu_pa_msg [CHECK_PARALLELISM-1:0];
ram_pageAlign_interface_partial_col_1_3_5_7_9 #(
	.QUAN_SIZE(QUAN_SIZE),
	.CHECK_PARALLELISM(CHECK_PARALLELISM),
	.LAYER_NUM(LAYER_NUM)
) vnu_ram_pageAlign_interface_submatrix_1_3_5_7_9 (
	.msg_out_0			(vnu_pa_msg[0]),
	.msg_out_1			(vnu_pa_msg[1]),
	.msg_out_2			(vnu_pa_msg[2]),
	.msg_out_3			(vnu_pa_msg[3]),
	.msg_out_4			(vnu_pa_msg[4]),
	.msg_out_5			(vnu_pa_msg[5]),
	.msg_out_6			(vnu_pa_msg[6]),
	.msg_out_7			(vnu_pa_msg[7]),
	.msg_out_8			(vnu_pa_msg[8]),
	.msg_out_9			(vnu_pa_msg[9]),
	.msg_out_10			(vnu_pa_msg[10]),
	.msg_out_11			(vnu_pa_msg[11]),
	.msg_out_12			(vnu_pa_msg[12]),
	.msg_out_13			(vnu_pa_msg[13]),
	.msg_out_14			(vnu_pa_msg[14]),
	.msg_out_15			(vnu_pa_msg[15]),
	.msg_out_16			(vnu_pa_msg[16]),
	.msg_out_17			(vnu_pa_msg[17]),
	.msg_out_18			(vnu_pa_msg[18]),
	.msg_out_19			(vnu_pa_msg[19]),
	.msg_out_20			(vnu_pa_msg[20]),
	.msg_out_21			(vnu_pa_msg[21]),
	.msg_out_22			(vnu_pa_msg[22]),
	.msg_out_23			(vnu_pa_msg[23]),
	.msg_out_24			(vnu_pa_msg[24]),
	.msg_out_25			(vnu_pa_msg[25]),
	.msg_out_26			(vnu_pa_msg[26]),
	.msg_out_27			(vnu_pa_msg[27]),
	.msg_out_28			(vnu_pa_msg[28]),
	.msg_out_29			(vnu_pa_msg[29]),
	.msg_out_30			(vnu_pa_msg[30]),
	.msg_out_31			(vnu_pa_msg[31]),
	.msg_out_32			(vnu_pa_msg[32]),
	.msg_out_33			(vnu_pa_msg[33]),
	.msg_out_34			(vnu_pa_msg[34]),
	.msg_out_35			(vnu_pa_msg[35]),
	.msg_out_36			(vnu_pa_msg[36]),
	.msg_out_37			(vnu_pa_msg[37]),
	.msg_out_38			(vnu_pa_msg[38]),
	.msg_out_39			(vnu_pa_msg[39]),
	.msg_out_40			(vnu_pa_msg[40]),
	.msg_out_41			(vnu_pa_msg[41]),
	.msg_out_42			(vnu_pa_msg[42]),
	.msg_out_43			(vnu_pa_msg[43]),
	.msg_out_44			(vnu_pa_msg[44]),
	.msg_out_45			(vnu_pa_msg[45]),
	.msg_out_46			(vnu_pa_msg[46]),
	.msg_out_47			(vnu_pa_msg[47]),
	.msg_out_48			(vnu_pa_msg[48]),
	.msg_out_49			(vnu_pa_msg[49]),
	.msg_out_50			(vnu_pa_msg[50]),
	.msg_out_51			(vnu_pa_msg[51]),
	.msg_out_52			(vnu_pa_msg[52]),
	.msg_out_53			(vnu_pa_msg[53]),
	.msg_out_54			(vnu_pa_msg[54]),
	.msg_out_55			(vnu_pa_msg[55]),
	.msg_out_56			(vnu_pa_msg[56]),
	.msg_out_57			(vnu_pa_msg[57]),
	.msg_out_58			(vnu_pa_msg[58]),
	.msg_out_59			(vnu_pa_msg[59]),
	.msg_out_60			(vnu_pa_msg[60]),
	.msg_out_61			(vnu_pa_msg[61]),
	.msg_out_62			(vnu_pa_msg[62]),
	.msg_out_63			(vnu_pa_msg[63]),
	.msg_out_64			(vnu_pa_msg[64]),
	.msg_out_65			(vnu_pa_msg[65]),
	.msg_out_66			(vnu_pa_msg[66]),
	.msg_out_67			(vnu_pa_msg[67]),
	.msg_out_68			(vnu_pa_msg[68]),
	.msg_out_69			(vnu_pa_msg[69]),
	.msg_out_70			(vnu_pa_msg[70]),
	.msg_out_71			(vnu_pa_msg[71]),
	.msg_out_72			(vnu_pa_msg[72]),
	.msg_out_73			(vnu_pa_msg[73]),
	.msg_out_74			(vnu_pa_msg[74]),
	.msg_out_75			(vnu_pa_msg[75]),
	.msg_out_76			(vnu_pa_msg[76]),
	.msg_out_77			(vnu_pa_msg[77]),
	.msg_out_78			(vnu_pa_msg[78]),
	.msg_out_79			(vnu_pa_msg[79]),
	.msg_out_80			(vnu_pa_msg[80]),
	.msg_out_81			(vnu_pa_msg[81]),
	.msg_out_82			(vnu_pa_msg[82]),
	.msg_out_83			(vnu_pa_msg[83]),
	.msg_out_84			(vnu_pa_msg[84]),
	.msg_out_85			(vnu_pa_msg[85]),
	.msg_out_86			(vnu_pa_msg[86]),
	.msg_out_87			(vnu_pa_msg[87]),
	.msg_out_88			(vnu_pa_msg[88]),
	.msg_out_89			(vnu_pa_msg[89]),
	.msg_out_90			(vnu_pa_msg[90]),
	.msg_out_91			(vnu_pa_msg[91]),
	.msg_out_92			(vnu_pa_msg[92]),
	.msg_out_93			(vnu_pa_msg[93]),
	.msg_out_94			(vnu_pa_msg[94]),
	.msg_out_95			(vnu_pa_msg[95]),
	.msg_out_96			(vnu_pa_msg[96]),
	.msg_out_97			(vnu_pa_msg[97]),
	.msg_out_98			(vnu_pa_msg[98]),
	.msg_out_99			(vnu_pa_msg[99]),
	.msg_out_100			(vnu_pa_msg[100]),
	.msg_out_101			(vnu_pa_msg[101]),
	.msg_out_102			(vnu_pa_msg[102]),
	.msg_out_103			(vnu_pa_msg[103]),
	.msg_out_104			(vnu_pa_msg[104]),
	.msg_out_105			(vnu_pa_msg[105]),
	.msg_out_106			(vnu_pa_msg[106]),
	.msg_out_107			(vnu_pa_msg[107]),
	.msg_out_108			(vnu_pa_msg[108]),
	.msg_out_109			(vnu_pa_msg[109]),
	.msg_out_110			(vnu_pa_msg[110]),
	.msg_out_111			(vnu_pa_msg[111]),
	.msg_out_112			(vnu_pa_msg[112]),
	.msg_out_113			(vnu_pa_msg[113]),
	.msg_out_114			(vnu_pa_msg[114]),
	.msg_out_115			(vnu_pa_msg[115]),
	.msg_out_116			(vnu_pa_msg[116]),
	.msg_out_117			(vnu_pa_msg[117]),
	.msg_out_118			(vnu_pa_msg[118]),
	.msg_out_119			(vnu_pa_msg[119]),
	.msg_out_120			(vnu_pa_msg[120]),
	.msg_out_121			(vnu_pa_msg[121]),
	.msg_out_122			(vnu_pa_msg[122]),
	.msg_out_123			(vnu_pa_msg[123]),
	.msg_out_124			(vnu_pa_msg[124]),
	.msg_out_125			(vnu_pa_msg[125]),
	.msg_out_126			(vnu_pa_msg[126]),
	.msg_out_127			(vnu_pa_msg[127]),
	.msg_out_128			(vnu_pa_msg[128]),
	.msg_out_129			(vnu_pa_msg[129]),
	.msg_out_130			(vnu_pa_msg[130]),
	.msg_out_131			(vnu_pa_msg[131]),
	.msg_out_132			(vnu_pa_msg[132]),
	.msg_out_133			(vnu_pa_msg[133]),
	.msg_out_134			(vnu_pa_msg[134]),
	.msg_out_135			(vnu_pa_msg[135]),
	.msg_out_136			(vnu_pa_msg[136]),
	.msg_out_137			(vnu_pa_msg[137]),
	.msg_out_138			(vnu_pa_msg[138]),
	.msg_out_139			(vnu_pa_msg[139]),
	.msg_out_140			(vnu_pa_msg[140]),
	.msg_out_141			(vnu_pa_msg[141]),
	.msg_out_142			(vnu_pa_msg[142]),
	.msg_out_143			(vnu_pa_msg[143]),
	.msg_out_144			(vnu_pa_msg[144]),
	.msg_out_145			(vnu_pa_msg[145]),
	.msg_out_146			(vnu_pa_msg[146]),
	.msg_out_147			(vnu_pa_msg[147]),
	.msg_out_148			(vnu_pa_msg[148]),
	.msg_out_149			(vnu_pa_msg[149]),
	.msg_out_150			(vnu_pa_msg[150]),
	.msg_out_151			(vnu_pa_msg[151]),
	.msg_out_152			(vnu_pa_msg[152]),
	.msg_out_153			(vnu_pa_msg[153]),
	.msg_out_154			(vnu_pa_msg[154]),
	.msg_out_155			(vnu_pa_msg[155]),
	.msg_out_156			(vnu_pa_msg[156]),
	.msg_out_157			(vnu_pa_msg[157]),
	.msg_out_158			(vnu_pa_msg[158]),
	.msg_out_159			(vnu_pa_msg[159]),
	.msg_out_160			(vnu_pa_msg[160]),
	.msg_out_161			(vnu_pa_msg[161]),
	.msg_out_162			(vnu_pa_msg[162]),
	.msg_out_163			(vnu_pa_msg[163]),
	.msg_out_164			(vnu_pa_msg[164]),
	.msg_out_165			(vnu_pa_msg[165]),
	.msg_out_166			(vnu_pa_msg[166]),
	.msg_out_167			(vnu_pa_msg[167]),
	.msg_out_168			(vnu_pa_msg[168]),
	.msg_out_169			(vnu_pa_msg[169]),
	.msg_out_170			(vnu_pa_msg[170]),
	.msg_out_171			(vnu_pa_msg[171]),
	.msg_out_172			(vnu_pa_msg[172]),
	.msg_out_173			(vnu_pa_msg[173]),
	.msg_out_174			(vnu_pa_msg[174]),
	.msg_out_175			(vnu_pa_msg[175]),
	.msg_out_176			(vnu_pa_msg[176]),
	.msg_out_177			(vnu_pa_msg[177]),
	.msg_out_178			(vnu_pa_msg[178]),
	.msg_out_179			(vnu_pa_msg[179]),
	.msg_out_180			(vnu_pa_msg[180]),
	.msg_out_181			(vnu_pa_msg[181]),
	.msg_out_182			(vnu_pa_msg[182]),
	.msg_out_183			(vnu_pa_msg[183]),
	.msg_out_184			(vnu_pa_msg[184]),
	.msg_out_185			(vnu_pa_msg[185]),
	.msg_out_186			(vnu_pa_msg[186]),
	.msg_out_187			(vnu_pa_msg[187]),
	.msg_out_188			(vnu_pa_msg[188]),
	.msg_out_189			(vnu_pa_msg[189]),
	.msg_out_190			(vnu_pa_msg[190]),
	.msg_out_191			(vnu_pa_msg[191]),
	.msg_out_192			(vnu_pa_msg[192]),
	.msg_out_193			(vnu_pa_msg[193]),
	.msg_out_194			(vnu_pa_msg[194]),
	.msg_out_195			(vnu_pa_msg[195]),
	.msg_out_196			(vnu_pa_msg[196]),
	.msg_out_197			(vnu_pa_msg[197]),
	.msg_out_198			(vnu_pa_msg[198]),
	.msg_out_199			(vnu_pa_msg[199]),
	.msg_out_200			(vnu_pa_msg[200]),
	.msg_out_201			(vnu_pa_msg[201]),
	.msg_out_202			(vnu_pa_msg[202]),
	.msg_out_203			(vnu_pa_msg[203]),
	.msg_out_204			(vnu_pa_msg[204]),
	.msg_out_205			(vnu_pa_msg[205]),
	.msg_out_206			(vnu_pa_msg[206]),
	.msg_out_207			(vnu_pa_msg[207]),
	.msg_out_208			(vnu_pa_msg[208]),
	.msg_out_209			(vnu_pa_msg[209]),
	.msg_out_210			(vnu_pa_msg[210]),
	.msg_out_211			(vnu_pa_msg[211]),
	.msg_out_212			(vnu_pa_msg[212]),
	.msg_out_213			(vnu_pa_msg[213]),
	.msg_out_214			(vnu_pa_msg[214]),
	.msg_out_215			(vnu_pa_msg[215]),
	.msg_out_216			(vnu_pa_msg[216]),
	.msg_out_217			(vnu_pa_msg[217]),
	.msg_out_218			(vnu_pa_msg[218]),
	.msg_out_219			(vnu_pa_msg[219]),
	.msg_out_220			(vnu_pa_msg[220]),
	.msg_out_221			(vnu_pa_msg[221]),
	.msg_out_222			(vnu_pa_msg[222]),
	.msg_out_223			(vnu_pa_msg[223]),
	.msg_out_224			(vnu_pa_msg[224]),
	.msg_out_225			(vnu_pa_msg[225]),
	.msg_out_226			(vnu_pa_msg[226]),
	.msg_out_227			(vnu_pa_msg[227]),
	.msg_out_228			(vnu_pa_msg[228]),
	.msg_out_229			(vnu_pa_msg[229]),
	.msg_out_230			(vnu_pa_msg[230]),
	.msg_out_231			(vnu_pa_msg[231]),
	.msg_out_232			(vnu_pa_msg[232]),
	.msg_out_233			(vnu_pa_msg[233]),
	.msg_out_234			(vnu_pa_msg[234]),
	.msg_out_235			(vnu_pa_msg[235]),
	.msg_out_236			(vnu_pa_msg[236]),
	.msg_out_237			(vnu_pa_msg[237]),
	.msg_out_238			(vnu_pa_msg[238]),
	.msg_out_239			(vnu_pa_msg[239]),
	.msg_out_240			(vnu_pa_msg[240]),
	.msg_out_241			(vnu_pa_msg[241]),
	.msg_out_242			(vnu_pa_msg[242]),
	.msg_out_243			(vnu_pa_msg[243]),
	.msg_out_244			(vnu_pa_msg[244]),
	.msg_out_245			(vnu_pa_msg[245]),
	.msg_out_246			(vnu_pa_msg[246]),
	.msg_out_247			(vnu_pa_msg[247]),
	.msg_out_248			(vnu_pa_msg[248]),
	.msg_out_249			(vnu_pa_msg[249]),
	.msg_out_250			(vnu_pa_msg[250]),
	.msg_out_251			(vnu_pa_msg[251]),
	.msg_out_252			(vnu_pa_msg[252]),
	.msg_out_253			(vnu_pa_msg[253]),
	.msg_out_254			(vnu_pa_msg[254]),
	.msg_in_0			(vnu_to_mem_0),
	.msg_in_1			(vnu_to_mem_1),
	.msg_in_2			(vnu_to_mem_2),
	.msg_in_3			(vnu_to_mem_3),
	.msg_in_4			(vnu_to_mem_4),
	.msg_in_5			(vnu_to_mem_5),
	.msg_in_6			(vnu_to_mem_6),
	.msg_in_7			(vnu_to_mem_7),
	.msg_in_8			(vnu_to_mem_8),
	.msg_in_9			(vnu_to_mem_9),
	.msg_in_10			(vnu_to_mem_10),
	.msg_in_11			(vnu_to_mem_11),
	.msg_in_12			(vnu_to_mem_12),
	.msg_in_13			(vnu_to_mem_13),
	.msg_in_14			(vnu_to_mem_14),
	.msg_in_15			(vnu_to_mem_15),
	.msg_in_16			(vnu_to_mem_16),
	.msg_in_17			(vnu_to_mem_17),
	.msg_in_18			(vnu_to_mem_18),
	.msg_in_19			(vnu_to_mem_19),
	.msg_in_20			(vnu_to_mem_20),
	.msg_in_21			(vnu_to_mem_21),
	.msg_in_22			(vnu_to_mem_22),
	.msg_in_23			(vnu_to_mem_23),
	.msg_in_24			(vnu_to_mem_24),
	.msg_in_25			(vnu_to_mem_25),
	.msg_in_26			(vnu_to_mem_26),
	.msg_in_27			(vnu_to_mem_27),
	.msg_in_28			(vnu_to_mem_28),
	.msg_in_29			(vnu_to_mem_29),
	.msg_in_30			(vnu_to_mem_30),
	.msg_in_31			(vnu_to_mem_31),
	.msg_in_32			(vnu_to_mem_32),
	.msg_in_33			(vnu_to_mem_33),
	.msg_in_34			(vnu_to_mem_34),
	.msg_in_35			(vnu_to_mem_35),
	.msg_in_36			(vnu_to_mem_36),
	.msg_in_37			(vnu_to_mem_37),
	.msg_in_38			(vnu_to_mem_38),
	.msg_in_39			(vnu_to_mem_39),
	.msg_in_40			(vnu_to_mem_40),
	.msg_in_41			(vnu_to_mem_41),
	.msg_in_42			(vnu_to_mem_42),
	.msg_in_43			(vnu_to_mem_43),
	.msg_in_44			(vnu_to_mem_44),
	.msg_in_45			(vnu_to_mem_45),
	.msg_in_46			(vnu_to_mem_46),
	.msg_in_47			(vnu_to_mem_47),
	.msg_in_48			(vnu_to_mem_48),
	.msg_in_49			(vnu_to_mem_49),
	.msg_in_50			(vnu_to_mem_50),
	.msg_in_51			(vnu_to_mem_51),
	.msg_in_52			(vnu_to_mem_52),
	.msg_in_53			(vnu_to_mem_53),
	.msg_in_54			(vnu_to_mem_54),
	.msg_in_55			(vnu_to_mem_55),
	.msg_in_56			(vnu_to_mem_56),
	.msg_in_57			(vnu_to_mem_57),
	.msg_in_58			(vnu_to_mem_58),
	.msg_in_59			(vnu_to_mem_59),
	.msg_in_60			(vnu_to_mem_60),
	.msg_in_61			(vnu_to_mem_61),
	.msg_in_62			(vnu_to_mem_62),
	.msg_in_63			(vnu_to_mem_63),
	.msg_in_64			(vnu_to_mem_64),
	.msg_in_65			(vnu_to_mem_65),
	.msg_in_66			(vnu_to_mem_66),
	.msg_in_67			(vnu_to_mem_67),
	.msg_in_68			(vnu_to_mem_68),
	.msg_in_69			(vnu_to_mem_69),
	.msg_in_70			(vnu_to_mem_70),
	.msg_in_71			(vnu_to_mem_71),
	.msg_in_72			(vnu_to_mem_72),
	.msg_in_73			(vnu_to_mem_73),
	.msg_in_74			(vnu_to_mem_74),
	.msg_in_75			(vnu_to_mem_75),
	.msg_in_76			(vnu_to_mem_76),
	.msg_in_77			(vnu_to_mem_77),
	.msg_in_78			(vnu_to_mem_78),
	.msg_in_79			(vnu_to_mem_79),
	.msg_in_80			(vnu_to_mem_80),
	.msg_in_81			(vnu_to_mem_81),
	.msg_in_82			(vnu_to_mem_82),
	.msg_in_83			(vnu_to_mem_83),
	.msg_in_84			(vnu_to_mem_84),
	.msg_in_85			(vnu_to_mem_85),
	.msg_in_86			(vnu_to_mem_86),
	.msg_in_87			(vnu_to_mem_87),
	.msg_in_88			(vnu_to_mem_88),
	.msg_in_89			(vnu_to_mem_89),
	.msg_in_90			(vnu_to_mem_90),
	.msg_in_91			(vnu_to_mem_91),
	.msg_in_92			(vnu_to_mem_92),
	.msg_in_93			(vnu_to_mem_93),
	.msg_in_94			(vnu_to_mem_94),
	.msg_in_95			(vnu_to_mem_95),
	.msg_in_96			(vnu_to_mem_96),
	.msg_in_97			(vnu_to_mem_97),
	.msg_in_98			(vnu_to_mem_98),
	.msg_in_99			(vnu_to_mem_99),
	.msg_in_100			(vnu_to_mem_100),
	.msg_in_101			(vnu_to_mem_101),
	.msg_in_102			(vnu_to_mem_102),
	.msg_in_103			(vnu_to_mem_103),
	.msg_in_104			(vnu_to_mem_104),
	.msg_in_105			(vnu_to_mem_105),
	.msg_in_106			(vnu_to_mem_106),
	.msg_in_107			(vnu_to_mem_107),
	.msg_in_108			(vnu_to_mem_108),
	.msg_in_109			(vnu_to_mem_109),
	.msg_in_110			(vnu_to_mem_110),
	.msg_in_111			(vnu_to_mem_111),
	.msg_in_112			(vnu_to_mem_112),
	.msg_in_113			(vnu_to_mem_113),
	.msg_in_114			(vnu_to_mem_114),
	.msg_in_115			(vnu_to_mem_115),
	.msg_in_116			(vnu_to_mem_116),
	.msg_in_117			(vnu_to_mem_117),
	.msg_in_118			(vnu_to_mem_118),
	.msg_in_119			(vnu_to_mem_119),
	.msg_in_120			(vnu_to_mem_120),
	.msg_in_121			(vnu_to_mem_121),
	.msg_in_122			(vnu_to_mem_122),
	.msg_in_123			(vnu_to_mem_123),
	.msg_in_124			(vnu_to_mem_124),
	.msg_in_125			(vnu_to_mem_125),
	.msg_in_126			(vnu_to_mem_126),
	.msg_in_127			(vnu_to_mem_127),
	.msg_in_128			(vnu_to_mem_128),
	.msg_in_129			(vnu_to_mem_129),
	.msg_in_130			(vnu_to_mem_130),
	.msg_in_131			(vnu_to_mem_131),
	.msg_in_132			(vnu_to_mem_132),
	.msg_in_133			(vnu_to_mem_133),
	.msg_in_134			(vnu_to_mem_134),
	.msg_in_135			(vnu_to_mem_135),
	.msg_in_136			(vnu_to_mem_136),
	.msg_in_137			(vnu_to_mem_137),
	.msg_in_138			(vnu_to_mem_138),
	.msg_in_139			(vnu_to_mem_139),
	.msg_in_140			(vnu_to_mem_140),
	.msg_in_141			(vnu_to_mem_141),
	.msg_in_142			(vnu_to_mem_142),
	.msg_in_143			(vnu_to_mem_143),
	.msg_in_144			(vnu_to_mem_144),
	.msg_in_145			(vnu_to_mem_145),
	.msg_in_146			(vnu_to_mem_146),
	.msg_in_147			(vnu_to_mem_147),
	.msg_in_148			(vnu_to_mem_148),
	.msg_in_149			(vnu_to_mem_149),
	.msg_in_150			(vnu_to_mem_150),
	.msg_in_151			(vnu_to_mem_151),
	.msg_in_152			(vnu_to_mem_152),
	.msg_in_153			(vnu_to_mem_153),
	.msg_in_154			(vnu_to_mem_154),
	.msg_in_155			(vnu_to_mem_155),
	.msg_in_156			(vnu_to_mem_156),
	.msg_in_157			(vnu_to_mem_157),
	.msg_in_158			(vnu_to_mem_158),
	.msg_in_159			(vnu_to_mem_159),
	.msg_in_160			(vnu_to_mem_160),
	.msg_in_161			(vnu_to_mem_161),
	.msg_in_162			(vnu_to_mem_162),
	.msg_in_163			(vnu_to_mem_163),
	.msg_in_164			(vnu_to_mem_164),
	.msg_in_165			(vnu_to_mem_165),
	.msg_in_166			(vnu_to_mem_166),
	.msg_in_167			(vnu_to_mem_167),
	.msg_in_168			(vnu_to_mem_168),
	.msg_in_169			(vnu_to_mem_169),
	.msg_in_170			(vnu_to_mem_170),
	.msg_in_171			(vnu_to_mem_171),
	.msg_in_172			(vnu_to_mem_172),
	.msg_in_173			(vnu_to_mem_173),
	.msg_in_174			(vnu_to_mem_174),
	.msg_in_175			(vnu_to_mem_175),
	.msg_in_176			(vnu_to_mem_176),
	.msg_in_177			(vnu_to_mem_177),
	.msg_in_178			(vnu_to_mem_178),
	.msg_in_179			(vnu_to_mem_179),
	.msg_in_180			(vnu_to_mem_180),
	.msg_in_181			(vnu_to_mem_181),
	.msg_in_182			(vnu_to_mem_182),
	.msg_in_183			(vnu_to_mem_183),
	.msg_in_184			(vnu_to_mem_184),
	.msg_in_185			(vnu_to_mem_185),
	.msg_in_186			(vnu_to_mem_186),
	.msg_in_187			(vnu_to_mem_187),
	.msg_in_188			(vnu_to_mem_188),
	.msg_in_189			(vnu_to_mem_189),
	.msg_in_190			(vnu_to_mem_190),
	.msg_in_191			(vnu_to_mem_191),
	.msg_in_192			(vnu_to_mem_192),
	.msg_in_193			(vnu_to_mem_193),
	.msg_in_194			(vnu_to_mem_194),
	.msg_in_195			(vnu_to_mem_195),
	.msg_in_196			(vnu_to_mem_196),
	.msg_in_197			(vnu_to_mem_197),
	.msg_in_198			(vnu_to_mem_198),
	.msg_in_199			(vnu_to_mem_199),
	.msg_in_200			(vnu_to_mem_200),
	.msg_in_201			(vnu_to_mem_201),
	.msg_in_202			(vnu_to_mem_202),
	.msg_in_203			(vnu_to_mem_203),
	.msg_in_204			(vnu_to_mem_204),
	.msg_in_205			(vnu_to_mem_205),
	.msg_in_206			(vnu_to_mem_206),
	.msg_in_207			(vnu_to_mem_207),
	.msg_in_208			(vnu_to_mem_208),
	.msg_in_209			(vnu_to_mem_209),
	.msg_in_210			(vnu_to_mem_210),
	.msg_in_211			(vnu_to_mem_211),
	.msg_in_212			(vnu_to_mem_212),
	.msg_in_213			(vnu_to_mem_213),
	.msg_in_214			(vnu_to_mem_214),
	.msg_in_215			(vnu_to_mem_215),
	.msg_in_216			(vnu_to_mem_216),
	.msg_in_217			(vnu_to_mem_217),
	.msg_in_218			(vnu_to_mem_218),
	.msg_in_219			(vnu_to_mem_219),
	.msg_in_220			(vnu_to_mem_220),
	.msg_in_221			(vnu_to_mem_221),
	.msg_in_222			(vnu_to_mem_222),
	.msg_in_223			(vnu_to_mem_223),
	.msg_in_224			(vnu_to_mem_224),
	.msg_in_225			(vnu_to_mem_225),
	.msg_in_226			(vnu_to_mem_226),
	.msg_in_227			(vnu_to_mem_227),
	.msg_in_228			(vnu_to_mem_228),
	.msg_in_229			(vnu_to_mem_229),
	.msg_in_230			(vnu_to_mem_230),
	.msg_in_231			(vnu_to_mem_231),
	.msg_in_232			(vnu_to_mem_232),
	.msg_in_233			(vnu_to_mem_233),
	.msg_in_234			(vnu_to_mem_234),
	.msg_in_235			(vnu_to_mem_235),
	.msg_in_236			(vnu_to_mem_236),
	.msg_in_237			(vnu_to_mem_237),
	.msg_in_238			(vnu_to_mem_238),
	.msg_in_239			(vnu_to_mem_239),
	.msg_in_240			(vnu_to_mem_240),
	.msg_in_241			(vnu_to_mem_241),
	.msg_in_242			(vnu_to_mem_242),
	.msg_in_243			(vnu_to_mem_243),
	.msg_in_244			(vnu_to_mem_244),
	.msg_in_245			(vnu_to_mem_245),
	.msg_in_246			(vnu_to_mem_246),
	.msg_in_247			(vnu_to_mem_247),
	.msg_in_248			(vnu_to_mem_248),
	.msg_in_249			(vnu_to_mem_249),
	.msg_in_250			(vnu_to_mem_250),
	.msg_in_251			(vnu_to_mem_251),
	.msg_in_252			(vnu_to_mem_252),
	.msg_in_253			(vnu_to_mem_253),
	.msg_in_254			(vnu_to_mem_254),
	.layer_status	(vnu_layer_status),
	.first_row_chunk	(last_row_chunk[1]),
	.sub_row_status	(vnu_sub_row_status[`ROW_SPLIT_FACTOR-1:0]),
	.sys_clk	(sys_clk),
	.rstn	(rstn)
);
/*-------------------------------------------------------*/
// Memory Instantiation
column_ram_pc255 #(
	.QUAN_SIZE(QUAN_SIZE),
	.CHECK_PARALLELISM(CHECK_PARALLELISM),
	.RAM_PORTA_RANGE(RAM_PORTA_RANGE),
	.RAM_PORTB_RANGE(RAM_PORTB_RANGE),
	.MEM_DEVICE_NUM(MEM_DEVICE_NUM),
	.DEPTH(DEPTH),
	.DATA_WIDTH(DATA_WIDTH),
	.FRAG_DATA_WIDTH(FRAG_DATA_WIDTH),
	.ADDR_WIDTH(ADDR_WIDTH)
) inst_column_ram_pc255 (
	.first_dout_0   (mem_to_cnu_0 ),
	.first_dout_1   (mem_to_cnu_1 ),
	.first_dout_2   (mem_to_cnu_2 ),
	.first_dout_3   (mem_to_cnu_3 ),
	.first_dout_4   (mem_to_cnu_4 ),
	.first_dout_5   (mem_to_cnu_5 ),
	.first_dout_6   (mem_to_cnu_6 ),
	.first_dout_7   (mem_to_cnu_7 ),
	.first_dout_8   (mem_to_cnu_8 ),
	.first_dout_9   (mem_to_cnu_9 ),
	.first_dout_10   (mem_to_cnu_10 ),
	.first_dout_11   (mem_to_cnu_11 ),
	.first_dout_12   (mem_to_cnu_12 ),
	.first_dout_13   (mem_to_cnu_13 ),
	.first_dout_14   (mem_to_cnu_14 ),
	.first_dout_15   (mem_to_cnu_15 ),
	.first_dout_16   (mem_to_cnu_16 ),
	.first_dout_17   (mem_to_cnu_17 ),
	.first_dout_18   (mem_to_cnu_18 ),
	.first_dout_19   (mem_to_cnu_19 ),
	.first_dout_20   (mem_to_cnu_20 ),
	.first_dout_21   (mem_to_cnu_21 ),
	.first_dout_22   (mem_to_cnu_22 ),
	.first_dout_23   (mem_to_cnu_23 ),
	.first_dout_24   (mem_to_cnu_24 ),
	.first_dout_25   (mem_to_cnu_25 ),
	.first_dout_26   (mem_to_cnu_26 ),
	.first_dout_27   (mem_to_cnu_27 ),
	.first_dout_28   (mem_to_cnu_28 ),
	.first_dout_29   (mem_to_cnu_29 ),
	.first_dout_30   (mem_to_cnu_30 ),
	.first_dout_31   (mem_to_cnu_31 ),
	.first_dout_32   (mem_to_cnu_32 ),
	.first_dout_33   (mem_to_cnu_33 ),
	.first_dout_34   (mem_to_cnu_34 ),
	.first_dout_35   (mem_to_cnu_35 ),
	.first_dout_36   (mem_to_cnu_36 ),
	.first_dout_37   (mem_to_cnu_37 ),
	.first_dout_38   (mem_to_cnu_38 ),
	.first_dout_39   (mem_to_cnu_39 ),
	.first_dout_40   (mem_to_cnu_40 ),
	.first_dout_41   (mem_to_cnu_41 ),
	.first_dout_42   (mem_to_cnu_42 ),
	.first_dout_43   (mem_to_cnu_43 ),
	.first_dout_44   (mem_to_cnu_44 ),
	.first_dout_45   (mem_to_cnu_45 ),
	.first_dout_46   (mem_to_cnu_46 ),
	.first_dout_47   (mem_to_cnu_47 ),
	.first_dout_48   (mem_to_cnu_48 ),
	.first_dout_49   (mem_to_cnu_49 ),
	.first_dout_50   (mem_to_cnu_50 ),
	.first_dout_51   (mem_to_cnu_51 ),
	.first_dout_52   (mem_to_cnu_52 ),
	.first_dout_53   (mem_to_cnu_53 ),
	.first_dout_54   (mem_to_cnu_54 ),
	.first_dout_55   (mem_to_cnu_55 ),
	.first_dout_56   (mem_to_cnu_56 ),
	.first_dout_57   (mem_to_cnu_57 ),
	.first_dout_58   (mem_to_cnu_58 ),
	.first_dout_59   (mem_to_cnu_59 ),
	.first_dout_60   (mem_to_cnu_60 ),
	.first_dout_61   (mem_to_cnu_61 ),
	.first_dout_62   (mem_to_cnu_62 ),
	.first_dout_63   (mem_to_cnu_63 ),
	.first_dout_64   (mem_to_cnu_64 ),
	.first_dout_65   (mem_to_cnu_65 ),
	.first_dout_66   (mem_to_cnu_66 ),
	.first_dout_67   (mem_to_cnu_67 ),
	.first_dout_68   (mem_to_cnu_68 ),
	.first_dout_69   (mem_to_cnu_69 ),
	.first_dout_70   (mem_to_cnu_70 ),
	.first_dout_71   (mem_to_cnu_71 ),
	.first_dout_72   (mem_to_cnu_72 ),
	.first_dout_73   (mem_to_cnu_73 ),
	.first_dout_74   (mem_to_cnu_74 ),
	.first_dout_75   (mem_to_cnu_75 ),
	.first_dout_76   (mem_to_cnu_76 ),
	.first_dout_77   (mem_to_cnu_77 ),
	.first_dout_78   (mem_to_cnu_78 ),
	.first_dout_79   (mem_to_cnu_79 ),
	.first_dout_80   (mem_to_cnu_80 ),
	.first_dout_81   (mem_to_cnu_81 ),
	.first_dout_82   (mem_to_cnu_82 ),
	.first_dout_83   (mem_to_cnu_83 ),
	.first_dout_84   (mem_to_cnu_84 ),
	.first_dout_85   (mem_to_cnu_85 ),
	.first_dout_86   (mem_to_cnu_86 ),
	.first_dout_87   (mem_to_cnu_87 ),
	.first_dout_88   (mem_to_cnu_88 ),
	.first_dout_89   (mem_to_cnu_89 ),
	.first_dout_90   (mem_to_cnu_90 ),
	.first_dout_91   (mem_to_cnu_91 ),
	.first_dout_92   (mem_to_cnu_92 ),
	.first_dout_93   (mem_to_cnu_93 ),
	.first_dout_94   (mem_to_cnu_94 ),
	.first_dout_95   (mem_to_cnu_95 ),
	.first_dout_96   (mem_to_cnu_96 ),
	.first_dout_97   (mem_to_cnu_97 ),
	.first_dout_98   (mem_to_cnu_98 ),
	.first_dout_99   (mem_to_cnu_99 ),
	.first_dout_100   (mem_to_cnu_100 ),
	.first_dout_101   (mem_to_cnu_101 ),
	.first_dout_102   (mem_to_cnu_102 ),
	.first_dout_103   (mem_to_cnu_103 ),
	.first_dout_104   (mem_to_cnu_104 ),
	.first_dout_105   (mem_to_cnu_105 ),
	.first_dout_106   (mem_to_cnu_106 ),
	.first_dout_107   (mem_to_cnu_107 ),
	.first_dout_108   (mem_to_cnu_108 ),
	.first_dout_109   (mem_to_cnu_109 ),
	.first_dout_110   (mem_to_cnu_110 ),
	.first_dout_111   (mem_to_cnu_111 ),
	.first_dout_112   (mem_to_cnu_112 ),
	.first_dout_113   (mem_to_cnu_113 ),
	.first_dout_114   (mem_to_cnu_114 ),
	.first_dout_115   (mem_to_cnu_115 ),
	.first_dout_116   (mem_to_cnu_116 ),
	.first_dout_117   (mem_to_cnu_117 ),
	.first_dout_118   (mem_to_cnu_118 ),
	.first_dout_119   (mem_to_cnu_119 ),
	.first_dout_120   (mem_to_cnu_120 ),
	.first_dout_121   (mem_to_cnu_121 ),
	.first_dout_122   (mem_to_cnu_122 ),
	.first_dout_123   (mem_to_cnu_123 ),
	.first_dout_124   (mem_to_cnu_124 ),
	.first_dout_125   (mem_to_cnu_125 ),
	.first_dout_126   (mem_to_cnu_126 ),
	.first_dout_127   (mem_to_cnu_127 ),
	.first_dout_128   (mem_to_cnu_128 ),
	.first_dout_129   (mem_to_cnu_129 ),
	.first_dout_130   (mem_to_cnu_130 ),
	.first_dout_131   (mem_to_cnu_131 ),
	.first_dout_132   (mem_to_cnu_132 ),
	.first_dout_133   (mem_to_cnu_133 ),
	.first_dout_134   (mem_to_cnu_134 ),
	.first_dout_135   (mem_to_cnu_135 ),
	.first_dout_136   (mem_to_cnu_136 ),
	.first_dout_137   (mem_to_cnu_137 ),
	.first_dout_138   (mem_to_cnu_138 ),
	.first_dout_139   (mem_to_cnu_139 ),
	.first_dout_140   (mem_to_cnu_140 ),
	.first_dout_141   (mem_to_cnu_141 ),
	.first_dout_142   (mem_to_cnu_142 ),
	.first_dout_143   (mem_to_cnu_143 ),
	.first_dout_144   (mem_to_cnu_144 ),
	.first_dout_145   (mem_to_cnu_145 ),
	.first_dout_146   (mem_to_cnu_146 ),
	.first_dout_147   (mem_to_cnu_147 ),
	.first_dout_148   (mem_to_cnu_148 ),
	.first_dout_149   (mem_to_cnu_149 ),
	.first_dout_150   (mem_to_cnu_150 ),
	.first_dout_151   (mem_to_cnu_151 ),
	.first_dout_152   (mem_to_cnu_152 ),
	.first_dout_153   (mem_to_cnu_153 ),
	.first_dout_154   (mem_to_cnu_154 ),
	.first_dout_155   (mem_to_cnu_155 ),
	.first_dout_156   (mem_to_cnu_156 ),
	.first_dout_157   (mem_to_cnu_157 ),
	.first_dout_158   (mem_to_cnu_158 ),
	.first_dout_159   (mem_to_cnu_159 ),
	.first_dout_160   (mem_to_cnu_160 ),
	.first_dout_161   (mem_to_cnu_161 ),
	.first_dout_162   (mem_to_cnu_162 ),
	.first_dout_163   (mem_to_cnu_163 ),
	.first_dout_164   (mem_to_cnu_164 ),
	.first_dout_165   (mem_to_cnu_165 ),
	.first_dout_166   (mem_to_cnu_166 ),
	.first_dout_167   (mem_to_cnu_167 ),
	.first_dout_168   (mem_to_cnu_168 ),
	.first_dout_169   (mem_to_cnu_169 ),
	.first_dout_170   (mem_to_cnu_170 ),
	.first_dout_171   (mem_to_cnu_171 ),
	.first_dout_172   (mem_to_cnu_172 ),
	.first_dout_173   (mem_to_cnu_173 ),
	.first_dout_174   (mem_to_cnu_174 ),
	.first_dout_175   (mem_to_cnu_175 ),
	.first_dout_176   (mem_to_cnu_176 ),
	.first_dout_177   (mem_to_cnu_177 ),
	.first_dout_178   (mem_to_cnu_178 ),
	.first_dout_179   (mem_to_cnu_179 ),
	.first_dout_180   (mem_to_cnu_180 ),
	.first_dout_181   (mem_to_cnu_181 ),
	.first_dout_182   (mem_to_cnu_182 ),
	.first_dout_183   (mem_to_cnu_183 ),
	.first_dout_184   (mem_to_cnu_184 ),
	.first_dout_185   (mem_to_cnu_185 ),
	.first_dout_186   (mem_to_cnu_186 ),
	.first_dout_187   (mem_to_cnu_187 ),
	.first_dout_188   (mem_to_cnu_188 ),
	.first_dout_189   (mem_to_cnu_189 ),
	.first_dout_190   (mem_to_cnu_190 ),
	.first_dout_191   (mem_to_cnu_191 ),
	.first_dout_192   (mem_to_cnu_192 ),
	.first_dout_193   (mem_to_cnu_193 ),
	.first_dout_194   (mem_to_cnu_194 ),
	.first_dout_195   (mem_to_cnu_195 ),
	.first_dout_196   (mem_to_cnu_196 ),
	.first_dout_197   (mem_to_cnu_197 ),
	.first_dout_198   (mem_to_cnu_198 ),
	.first_dout_199   (mem_to_cnu_199 ),
	.first_dout_200   (mem_to_cnu_200 ),
	.first_dout_201   (mem_to_cnu_201 ),
	.first_dout_202   (mem_to_cnu_202 ),
	.first_dout_203   (mem_to_cnu_203 ),
	.first_dout_204   (mem_to_cnu_204 ),
	.first_dout_205   (mem_to_cnu_205 ),
	.first_dout_206   (mem_to_cnu_206 ),
	.first_dout_207   (mem_to_cnu_207 ),
	.first_dout_208   (mem_to_cnu_208 ),
	.first_dout_209   (mem_to_cnu_209 ),
	.first_dout_210   (mem_to_cnu_210 ),
	.first_dout_211   (mem_to_cnu_211 ),
	.first_dout_212   (mem_to_cnu_212 ),
	.first_dout_213   (mem_to_cnu_213 ),
	.first_dout_214   (mem_to_cnu_214 ),
	.first_dout_215   (mem_to_cnu_215 ),
	.first_dout_216   (mem_to_cnu_216 ),
	.first_dout_217   (mem_to_cnu_217 ),
	.first_dout_218   (mem_to_cnu_218 ),
	.first_dout_219   (mem_to_cnu_219 ),
	.first_dout_220   (mem_to_cnu_220 ),
	.first_dout_221   (mem_to_cnu_221 ),
	.first_dout_222   (mem_to_cnu_222 ),
	.first_dout_223   (mem_to_cnu_223 ),
	.first_dout_224   (mem_to_cnu_224 ),
	.first_dout_225   (mem_to_cnu_225 ),
	.first_dout_226   (mem_to_cnu_226 ),
	.first_dout_227   (mem_to_cnu_227 ),
	.first_dout_228   (mem_to_cnu_228 ),
	.first_dout_229   (mem_to_cnu_229 ),
	.first_dout_230   (mem_to_cnu_230 ),
	.first_dout_231   (mem_to_cnu_231 ),
	.first_dout_232   (mem_to_cnu_232 ),
	.first_dout_233   (mem_to_cnu_233 ),
	.first_dout_234   (mem_to_cnu_234 ),
	.first_dout_235   (mem_to_cnu_235 ),
	.first_dout_236   (mem_to_cnu_236 ),
	.first_dout_237   (mem_to_cnu_237 ),
	.first_dout_238   (mem_to_cnu_238 ),
	.first_dout_239   (mem_to_cnu_239 ),
	.first_dout_240   (mem_to_cnu_240 ),
	.first_dout_241   (mem_to_cnu_241 ),
	.first_dout_242   (mem_to_cnu_242 ),
	.first_dout_243   (mem_to_cnu_243 ),
	.first_dout_244   (mem_to_cnu_244 ),
	.first_dout_245   (mem_to_cnu_245 ),
	.first_dout_246   (mem_to_cnu_246 ),
	.first_dout_247   (mem_to_cnu_247 ),
	.first_dout_248   (mem_to_cnu_248 ),
	.first_dout_249   (mem_to_cnu_249 ),
	.first_dout_250   (mem_to_cnu_250 ),
	.first_dout_251   (mem_to_cnu_251 ),
	.first_dout_252   (mem_to_cnu_252 ),
	.first_dout_253   (mem_to_cnu_253 ),
	.first_dout_254   (mem_to_cnu_254 ),

	.first_dout_0   (mem_to_cnu_0 ),
	.first_dout_1   (mem_to_cnu_1 ),
	.first_dout_2   (mem_to_cnu_2 ),
	.first_dout_3   (mem_to_cnu_3 ),
	.first_dout_4   (mem_to_cnu_4 ),
	.first_dout_5   (mem_to_cnu_5 ),
	.first_dout_6   (mem_to_cnu_6 ),
	.first_dout_7   (mem_to_cnu_7 ),
	.first_dout_8   (mem_to_cnu_8 ),
	.first_dout_9   (mem_to_cnu_9 ),
	.first_dout_10   (mem_to_cnu_10 ),
	.first_dout_11   (mem_to_cnu_11 ),
	.first_dout_12   (mem_to_cnu_12 ),
	.first_dout_13   (mem_to_cnu_13 ),
	.first_dout_14   (mem_to_cnu_14 ),
	.first_dout_15   (mem_to_cnu_15 ),
	.first_dout_16   (mem_to_cnu_16 ),
	.first_dout_17   (mem_to_cnu_17 ),
	.first_dout_18   (mem_to_cnu_18 ),
	.first_dout_19   (mem_to_cnu_19 ),
	.first_dout_20   (mem_to_cnu_20 ),
	.first_dout_21   (mem_to_cnu_21 ),
	.first_dout_22   (mem_to_cnu_22 ),
	.first_dout_23   (mem_to_cnu_23 ),
	.first_dout_24   (mem_to_cnu_24 ),
	.first_dout_25   (mem_to_cnu_25 ),
	.first_dout_26   (mem_to_cnu_26 ),
	.first_dout_27   (mem_to_cnu_27 ),
	.first_dout_28   (mem_to_cnu_28 ),
	.first_dout_29   (mem_to_cnu_29 ),
	.first_dout_30   (mem_to_cnu_30 ),
	.first_dout_31   (mem_to_cnu_31 ),
	.first_dout_32   (mem_to_cnu_32 ),
	.first_dout_33   (mem_to_cnu_33 ),
	.first_dout_34   (mem_to_cnu_34 ),
	.first_dout_35   (mem_to_cnu_35 ),
	.first_dout_36   (mem_to_cnu_36 ),
	.first_dout_37   (mem_to_cnu_37 ),
	.first_dout_38   (mem_to_cnu_38 ),
	.first_dout_39   (mem_to_cnu_39 ),
	.first_dout_40   (mem_to_cnu_40 ),
	.first_dout_41   (mem_to_cnu_41 ),
	.first_dout_42   (mem_to_cnu_42 ),
	.first_dout_43   (mem_to_cnu_43 ),
	.first_dout_44   (mem_to_cnu_44 ),
	.first_dout_45   (mem_to_cnu_45 ),
	.first_dout_46   (mem_to_cnu_46 ),
	.first_dout_47   (mem_to_cnu_47 ),
	.first_dout_48   (mem_to_cnu_48 ),
	.first_dout_49   (mem_to_cnu_49 ),
	.first_dout_50   (mem_to_cnu_50 ),
	.first_dout_51   (mem_to_cnu_51 ),
	.first_dout_52   (mem_to_cnu_52 ),
	.first_dout_53   (mem_to_cnu_53 ),
	.first_dout_54   (mem_to_cnu_54 ),
	.first_dout_55   (mem_to_cnu_55 ),
	.first_dout_56   (mem_to_cnu_56 ),
	.first_dout_57   (mem_to_cnu_57 ),
	.first_dout_58   (mem_to_cnu_58 ),
	.first_dout_59   (mem_to_cnu_59 ),
	.first_dout_60   (mem_to_cnu_60 ),
	.first_dout_61   (mem_to_cnu_61 ),
	.first_dout_62   (mem_to_cnu_62 ),
	.first_dout_63   (mem_to_cnu_63 ),
	.first_dout_64   (mem_to_cnu_64 ),
	.first_dout_65   (mem_to_cnu_65 ),
	.first_dout_66   (mem_to_cnu_66 ),
	.first_dout_67   (mem_to_cnu_67 ),
	.first_dout_68   (mem_to_cnu_68 ),
	.first_dout_69   (mem_to_cnu_69 ),
	.first_dout_70   (mem_to_cnu_70 ),
	.first_dout_71   (mem_to_cnu_71 ),
	.first_dout_72   (mem_to_cnu_72 ),
	.first_dout_73   (mem_to_cnu_73 ),
	.first_dout_74   (mem_to_cnu_74 ),
	.first_dout_75   (mem_to_cnu_75 ),
	.first_dout_76   (mem_to_cnu_76 ),
	.first_dout_77   (mem_to_cnu_77 ),
	.first_dout_78   (mem_to_cnu_78 ),
	.first_dout_79   (mem_to_cnu_79 ),
	.first_dout_80   (mem_to_cnu_80 ),
	.first_dout_81   (mem_to_cnu_81 ),
	.first_dout_82   (mem_to_cnu_82 ),
	.first_dout_83   (mem_to_cnu_83 ),
	.first_dout_84   (mem_to_cnu_84 ),
	.first_dout_85   (mem_to_cnu_85 ),
	.first_dout_86   (mem_to_cnu_86 ),
	.first_dout_87   (mem_to_cnu_87 ),
	.first_dout_88   (mem_to_cnu_88 ),
	.first_dout_89   (mem_to_cnu_89 ),
	.first_dout_90   (mem_to_cnu_90 ),
	.first_dout_91   (mem_to_cnu_91 ),
	.first_dout_92   (mem_to_cnu_92 ),
	.first_dout_93   (mem_to_cnu_93 ),
	.first_dout_94   (mem_to_cnu_94 ),
	.first_dout_95   (mem_to_cnu_95 ),
	.first_dout_96   (mem_to_cnu_96 ),
	.first_dout_97   (mem_to_cnu_97 ),
	.first_dout_98   (mem_to_cnu_98 ),
	.first_dout_99   (mem_to_cnu_99 ),
	.first_dout_100   (mem_to_cnu_100 ),
	.first_dout_101   (mem_to_cnu_101 ),
	.first_dout_102   (mem_to_cnu_102 ),
	.first_dout_103   (mem_to_cnu_103 ),
	.first_dout_104   (mem_to_cnu_104 ),
	.first_dout_105   (mem_to_cnu_105 ),
	.first_dout_106   (mem_to_cnu_106 ),
	.first_dout_107   (mem_to_cnu_107 ),
	.first_dout_108   (mem_to_cnu_108 ),
	.first_dout_109   (mem_to_cnu_109 ),
	.first_dout_110   (mem_to_cnu_110 ),
	.first_dout_111   (mem_to_cnu_111 ),
	.first_dout_112   (mem_to_cnu_112 ),
	.first_dout_113   (mem_to_cnu_113 ),
	.first_dout_114   (mem_to_cnu_114 ),
	.first_dout_115   (mem_to_cnu_115 ),
	.first_dout_116   (mem_to_cnu_116 ),
	.first_dout_117   (mem_to_cnu_117 ),
	.first_dout_118   (mem_to_cnu_118 ),
	.first_dout_119   (mem_to_cnu_119 ),
	.first_dout_120   (mem_to_cnu_120 ),
	.first_dout_121   (mem_to_cnu_121 ),
	.first_dout_122   (mem_to_cnu_122 ),
	.first_dout_123   (mem_to_cnu_123 ),
	.first_dout_124   (mem_to_cnu_124 ),
	.first_dout_125   (mem_to_cnu_125 ),
	.first_dout_126   (mem_to_cnu_126 ),
	.first_dout_127   (mem_to_cnu_127 ),
	.first_dout_128   (mem_to_cnu_128 ),
	.first_dout_129   (mem_to_cnu_129 ),
	.first_dout_130   (mem_to_cnu_130 ),
	.first_dout_131   (mem_to_cnu_131 ),
	.first_dout_132   (mem_to_cnu_132 ),
	.first_dout_133   (mem_to_cnu_133 ),
	.first_dout_134   (mem_to_cnu_134 ),
	.first_dout_135   (mem_to_cnu_135 ),
	.first_dout_136   (mem_to_cnu_136 ),
	.first_dout_137   (mem_to_cnu_137 ),
	.first_dout_138   (mem_to_cnu_138 ),
	.first_dout_139   (mem_to_cnu_139 ),
	.first_dout_140   (mem_to_cnu_140 ),
	.first_dout_141   (mem_to_cnu_141 ),
	.first_dout_142   (mem_to_cnu_142 ),
	.first_dout_143   (mem_to_cnu_143 ),
	.first_dout_144   (mem_to_cnu_144 ),
	.first_dout_145   (mem_to_cnu_145 ),
	.first_dout_146   (mem_to_cnu_146 ),
	.first_dout_147   (mem_to_cnu_147 ),
	.first_dout_148   (mem_to_cnu_148 ),
	.first_dout_149   (mem_to_cnu_149 ),
	.first_dout_150   (mem_to_cnu_150 ),
	.first_dout_151   (mem_to_cnu_151 ),
	.first_dout_152   (mem_to_cnu_152 ),
	.first_dout_153   (mem_to_cnu_153 ),
	.first_dout_154   (mem_to_cnu_154 ),
	.first_dout_155   (mem_to_cnu_155 ),
	.first_dout_156   (mem_to_cnu_156 ),
	.first_dout_157   (mem_to_cnu_157 ),
	.first_dout_158   (mem_to_cnu_158 ),
	.first_dout_159   (mem_to_cnu_159 ),
	.first_dout_160   (mem_to_cnu_160 ),
	.first_dout_161   (mem_to_cnu_161 ),
	.first_dout_162   (mem_to_cnu_162 ),
	.first_dout_163   (mem_to_cnu_163 ),
	.first_dout_164   (mem_to_cnu_164 ),
	.first_dout_165   (mem_to_cnu_165 ),
	.first_dout_166   (mem_to_cnu_166 ),
	.first_dout_167   (mem_to_cnu_167 ),
	.first_dout_168   (mem_to_cnu_168 ),
	.first_dout_169   (mem_to_cnu_169 ),
	.first_dout_170   (mem_to_cnu_170 ),
	.first_dout_171   (mem_to_cnu_171 ),
	.first_dout_172   (mem_to_cnu_172 ),
	.first_dout_173   (mem_to_cnu_173 ),
	.first_dout_174   (mem_to_cnu_174 ),
	.first_dout_175   (mem_to_cnu_175 ),
	.first_dout_176   (mem_to_cnu_176 ),
	.first_dout_177   (mem_to_cnu_177 ),
	.first_dout_178   (mem_to_cnu_178 ),
	.first_dout_179   (mem_to_cnu_179 ),
	.first_dout_180   (mem_to_cnu_180 ),
	.first_dout_181   (mem_to_cnu_181 ),
	.first_dout_182   (mem_to_cnu_182 ),
	.first_dout_183   (mem_to_cnu_183 ),
	.first_dout_184   (mem_to_cnu_184 ),
	.first_dout_185   (mem_to_cnu_185 ),
	.first_dout_186   (mem_to_cnu_186 ),
	.first_dout_187   (mem_to_cnu_187 ),
	.first_dout_188   (mem_to_cnu_188 ),
	.first_dout_189   (mem_to_cnu_189 ),
	.first_dout_190   (mem_to_cnu_190 ),
	.first_dout_191   (mem_to_cnu_191 ),
	.first_dout_192   (mem_to_cnu_192 ),
	.first_dout_193   (mem_to_cnu_193 ),
	.first_dout_194   (mem_to_cnu_194 ),
	.first_dout_195   (mem_to_cnu_195 ),
	.first_dout_196   (mem_to_cnu_196 ),
	.first_dout_197   (mem_to_cnu_197 ),
	.first_dout_198   (mem_to_cnu_198 ),
	.first_dout_199   (mem_to_cnu_199 ),
	.first_dout_200   (mem_to_cnu_200 ),
	.first_dout_201   (mem_to_cnu_201 ),
	.first_dout_202   (mem_to_cnu_202 ),
	.first_dout_203   (mem_to_cnu_203 ),
	.first_dout_204   (mem_to_cnu_204 ),
	.first_dout_205   (mem_to_cnu_205 ),
	.first_dout_206   (mem_to_cnu_206 ),
	.first_dout_207   (mem_to_cnu_207 ),
	.first_dout_208   (mem_to_cnu_208 ),
	.first_dout_209   (mem_to_cnu_209 ),
	.first_dout_210   (mem_to_cnu_210 ),
	.first_dout_211   (mem_to_cnu_211 ),
	.first_dout_212   (mem_to_cnu_212 ),
	.first_dout_213   (mem_to_cnu_213 ),
	.first_dout_214   (mem_to_cnu_214 ),
	.first_dout_215   (mem_to_cnu_215 ),
	.first_dout_216   (mem_to_cnu_216 ),
	.first_dout_217   (mem_to_cnu_217 ),
	.first_dout_218   (mem_to_cnu_218 ),
	.first_dout_219   (mem_to_cnu_219 ),
	.first_dout_220   (mem_to_cnu_220 ),
	.first_dout_221   (mem_to_cnu_221 ),
	.first_dout_222   (mem_to_cnu_222 ),
	.first_dout_223   (mem_to_cnu_223 ),
	.first_dout_224   (mem_to_cnu_224 ),
	.first_dout_225   (mem_to_cnu_225 ),
	.first_dout_226   (mem_to_cnu_226 ),
	.first_dout_227   (mem_to_cnu_227 ),
	.first_dout_228   (mem_to_cnu_228 ),
	.first_dout_229   (mem_to_cnu_229 ),
	.first_dout_230   (mem_to_cnu_230 ),
	.first_dout_231   (mem_to_cnu_231 ),
	.first_dout_232   (mem_to_cnu_232 ),
	.first_dout_233   (mem_to_cnu_233 ),
	.first_dout_234   (mem_to_cnu_234 ),
	.first_dout_235   (mem_to_cnu_235 ),
	.first_dout_236   (mem_to_cnu_236 ),
	.first_dout_237   (mem_to_cnu_237 ),
	.first_dout_238   (mem_to_cnu_238 ),
	.first_dout_239   (mem_to_cnu_239 ),
	.first_dout_240   (mem_to_cnu_240 ),
	.first_dout_241   (mem_to_cnu_241 ),
	.first_dout_242   (mem_to_cnu_242 ),
	.first_dout_243   (mem_to_cnu_243 ),
	.first_dout_244   (mem_to_cnu_244 ),
	.first_dout_245   (mem_to_cnu_245 ),
	.first_dout_246   (mem_to_cnu_246 ),
	.first_dout_247   (mem_to_cnu_247 ),
	.first_dout_248   (mem_to_cnu_248 ),
	.first_dout_249   (mem_to_cnu_249 ),
	.first_dout_250   (mem_to_cnu_250 ),
	.first_dout_251   (mem_to_cnu_251 ),
	.first_dout_252   (mem_to_cnu_252 ),
	.first_dout_253   (mem_to_cnu_253 ),
	.first_dout_254   (mem_to_cnu_254 ),

	.first_din_0    (cnu_pa_msg[0]),
	.first_din_1    (cnu_pa_msg[1]),
	.first_din_2    (cnu_pa_msg[2]),
	.first_din_3    (cnu_pa_msg[3]),
	.first_din_4    (cnu_pa_msg[4]),
	.first_din_5    (cnu_pa_msg[5]),
	.first_din_6    (cnu_pa_msg[6]),
	.first_din_7    (cnu_pa_msg[7]),
	.first_din_8    (cnu_pa_msg[8]),
	.first_din_9    (cnu_pa_msg[9]),
	.first_din_10    (cnu_pa_msg[10]),
	.first_din_11    (cnu_pa_msg[11]),
	.first_din_12    (cnu_pa_msg[12]),
	.first_din_13    (cnu_pa_msg[13]),
	.first_din_14    (cnu_pa_msg[14]),
	.first_din_15    (cnu_pa_msg[15]),
	.first_din_16    (cnu_pa_msg[16]),
	.first_din_17    (cnu_pa_msg[17]),
	.first_din_18    (cnu_pa_msg[18]),
	.first_din_19    (cnu_pa_msg[19]),
	.first_din_20    (cnu_pa_msg[20]),
	.first_din_21    (cnu_pa_msg[21]),
	.first_din_22    (cnu_pa_msg[22]),
	.first_din_23    (cnu_pa_msg[23]),
	.first_din_24    (cnu_pa_msg[24]),
	.first_din_25    (cnu_pa_msg[25]),
	.first_din_26    (cnu_pa_msg[26]),
	.first_din_27    (cnu_pa_msg[27]),
	.first_din_28    (cnu_pa_msg[28]),
	.first_din_29    (cnu_pa_msg[29]),
	.first_din_30    (cnu_pa_msg[30]),
	.first_din_31    (cnu_pa_msg[31]),
	.first_din_32    (cnu_pa_msg[32]),
	.first_din_33    (cnu_pa_msg[33]),
	.first_din_34    (cnu_pa_msg[34]),
	.first_din_35    (cnu_pa_msg[35]),
	.first_din_36    (cnu_pa_msg[36]),
	.first_din_37    (cnu_pa_msg[37]),
	.first_din_38    (cnu_pa_msg[38]),
	.first_din_39    (cnu_pa_msg[39]),
	.first_din_40    (cnu_pa_msg[40]),
	.first_din_41    (cnu_pa_msg[41]),
	.first_din_42    (cnu_pa_msg[42]),
	.first_din_43    (cnu_pa_msg[43]),
	.first_din_44    (cnu_pa_msg[44]),
	.first_din_45    (cnu_pa_msg[45]),
	.first_din_46    (cnu_pa_msg[46]),
	.first_din_47    (cnu_pa_msg[47]),
	.first_din_48    (cnu_pa_msg[48]),
	.first_din_49    (cnu_pa_msg[49]),
	.first_din_50    (cnu_pa_msg[50]),
	.first_din_51    (cnu_pa_msg[51]),
	.first_din_52    (cnu_pa_msg[52]),
	.first_din_53    (cnu_pa_msg[53]),
	.first_din_54    (cnu_pa_msg[54]),
	.first_din_55    (cnu_pa_msg[55]),
	.first_din_56    (cnu_pa_msg[56]),
	.first_din_57    (cnu_pa_msg[57]),
	.first_din_58    (cnu_pa_msg[58]),
	.first_din_59    (cnu_pa_msg[59]),
	.first_din_60    (cnu_pa_msg[60]),
	.first_din_61    (cnu_pa_msg[61]),
	.first_din_62    (cnu_pa_msg[62]),
	.first_din_63    (cnu_pa_msg[63]),
	.first_din_64    (cnu_pa_msg[64]),
	.first_din_65    (cnu_pa_msg[65]),
	.first_din_66    (cnu_pa_msg[66]),
	.first_din_67    (cnu_pa_msg[67]),
	.first_din_68    (cnu_pa_msg[68]),
	.first_din_69    (cnu_pa_msg[69]),
	.first_din_70    (cnu_pa_msg[70]),
	.first_din_71    (cnu_pa_msg[71]),
	.first_din_72    (cnu_pa_msg[72]),
	.first_din_73    (cnu_pa_msg[73]),
	.first_din_74    (cnu_pa_msg[74]),
	.first_din_75    (cnu_pa_msg[75]),
	.first_din_76    (cnu_pa_msg[76]),
	.first_din_77    (cnu_pa_msg[77]),
	.first_din_78    (cnu_pa_msg[78]),
	.first_din_79    (cnu_pa_msg[79]),
	.first_din_80    (cnu_pa_msg[80]),
	.first_din_81    (cnu_pa_msg[81]),
	.first_din_82    (cnu_pa_msg[82]),
	.first_din_83    (cnu_pa_msg[83]),
	.first_din_84    (cnu_pa_msg[84]),
	.first_din_85    (cnu_pa_msg[85]),
	.first_din_86    (cnu_pa_msg[86]),
	.first_din_87    (cnu_pa_msg[87]),
	.first_din_88    (cnu_pa_msg[88]),
	.first_din_89    (cnu_pa_msg[89]),
	.first_din_90    (cnu_pa_msg[90]),
	.first_din_91    (cnu_pa_msg[91]),
	.first_din_92    (cnu_pa_msg[92]),
	.first_din_93    (cnu_pa_msg[93]),
	.first_din_94    (cnu_pa_msg[94]),
	.first_din_95    (cnu_pa_msg[95]),
	.first_din_96    (cnu_pa_msg[96]),
	.first_din_97    (cnu_pa_msg[97]),
	.first_din_98    (cnu_pa_msg[98]),
	.first_din_99    (cnu_pa_msg[99]),
	.first_din_100    (cnu_pa_msg[100]),
	.first_din_101    (cnu_pa_msg[101]),
	.first_din_102    (cnu_pa_msg[102]),
	.first_din_103    (cnu_pa_msg[103]),
	.first_din_104    (cnu_pa_msg[104]),
	.first_din_105    (cnu_pa_msg[105]),
	.first_din_106    (cnu_pa_msg[106]),
	.first_din_107    (cnu_pa_msg[107]),
	.first_din_108    (cnu_pa_msg[108]),
	.first_din_109    (cnu_pa_msg[109]),
	.first_din_110    (cnu_pa_msg[110]),
	.first_din_111    (cnu_pa_msg[111]),
	.first_din_112    (cnu_pa_msg[112]),
	.first_din_113    (cnu_pa_msg[113]),
	.first_din_114    (cnu_pa_msg[114]),
	.first_din_115    (cnu_pa_msg[115]),
	.first_din_116    (cnu_pa_msg[116]),
	.first_din_117    (cnu_pa_msg[117]),
	.first_din_118    (cnu_pa_msg[118]),
	.first_din_119    (cnu_pa_msg[119]),
	.first_din_120    (cnu_pa_msg[120]),
	.first_din_121    (cnu_pa_msg[121]),
	.first_din_122    (cnu_pa_msg[122]),
	.first_din_123    (cnu_pa_msg[123]),
	.first_din_124    (cnu_pa_msg[124]),
	.first_din_125    (cnu_pa_msg[125]),
	.first_din_126    (cnu_pa_msg[126]),
	.first_din_127    (cnu_pa_msg[127]),
	.first_din_128    (cnu_pa_msg[128]),
	.first_din_129    (cnu_pa_msg[129]),
	.first_din_130    (cnu_pa_msg[130]),
	.first_din_131    (cnu_pa_msg[131]),
	.first_din_132    (cnu_pa_msg[132]),
	.first_din_133    (cnu_pa_msg[133]),
	.first_din_134    (cnu_pa_msg[134]),
	.first_din_135    (cnu_pa_msg[135]),
	.first_din_136    (cnu_pa_msg[136]),
	.first_din_137    (cnu_pa_msg[137]),
	.first_din_138    (cnu_pa_msg[138]),
	.first_din_139    (cnu_pa_msg[139]),
	.first_din_140    (cnu_pa_msg[140]),
	.first_din_141    (cnu_pa_msg[141]),
	.first_din_142    (cnu_pa_msg[142]),
	.first_din_143    (cnu_pa_msg[143]),
	.first_din_144    (cnu_pa_msg[144]),
	.first_din_145    (cnu_pa_msg[145]),
	.first_din_146    (cnu_pa_msg[146]),
	.first_din_147    (cnu_pa_msg[147]),
	.first_din_148    (cnu_pa_msg[148]),
	.first_din_149    (cnu_pa_msg[149]),
	.first_din_150    (cnu_pa_msg[150]),
	.first_din_151    (cnu_pa_msg[151]),
	.first_din_152    (cnu_pa_msg[152]),
	.first_din_153    (cnu_pa_msg[153]),
	.first_din_154    (cnu_pa_msg[154]),
	.first_din_155    (cnu_pa_msg[155]),
	.first_din_156    (cnu_pa_msg[156]),
	.first_din_157    (cnu_pa_msg[157]),
	.first_din_158    (cnu_pa_msg[158]),
	.first_din_159    (cnu_pa_msg[159]),
	.first_din_160    (cnu_pa_msg[160]),
	.first_din_161    (cnu_pa_msg[161]),
	.first_din_162    (cnu_pa_msg[162]),
	.first_din_163    (cnu_pa_msg[163]),
	.first_din_164    (cnu_pa_msg[164]),
	.first_din_165    (cnu_pa_msg[165]),
	.first_din_166    (cnu_pa_msg[166]),
	.first_din_167    (cnu_pa_msg[167]),
	.first_din_168    (cnu_pa_msg[168]),
	.first_din_169    (cnu_pa_msg[169]),
	.first_din_170    (cnu_pa_msg[170]),
	.first_din_171    (cnu_pa_msg[171]),
	.first_din_172    (cnu_pa_msg[172]),
	.first_din_173    (cnu_pa_msg[173]),
	.first_din_174    (cnu_pa_msg[174]),
	.first_din_175    (cnu_pa_msg[175]),
	.first_din_176    (cnu_pa_msg[176]),
	.first_din_177    (cnu_pa_msg[177]),
	.first_din_178    (cnu_pa_msg[178]),
	.first_din_179    (cnu_pa_msg[179]),
	.first_din_180    (cnu_pa_msg[180]),
	.first_din_181    (cnu_pa_msg[181]),
	.first_din_182    (cnu_pa_msg[182]),
	.first_din_183    (cnu_pa_msg[183]),
	.first_din_184    (cnu_pa_msg[184]),
	.first_din_185    (cnu_pa_msg[185]),
	.first_din_186    (cnu_pa_msg[186]),
	.first_din_187    (cnu_pa_msg[187]),
	.first_din_188    (cnu_pa_msg[188]),
	.first_din_189    (cnu_pa_msg[189]),
	.first_din_190    (cnu_pa_msg[190]),
	.first_din_191    (cnu_pa_msg[191]),
	.first_din_192    (cnu_pa_msg[192]),
	.first_din_193    (cnu_pa_msg[193]),
	.first_din_194    (cnu_pa_msg[194]),
	.first_din_195    (cnu_pa_msg[195]),
	.first_din_196    (cnu_pa_msg[196]),
	.first_din_197    (cnu_pa_msg[197]),
	.first_din_198    (cnu_pa_msg[198]),
	.first_din_199    (cnu_pa_msg[199]),
	.first_din_200    (cnu_pa_msg[200]),
	.first_din_201    (cnu_pa_msg[201]),
	.first_din_202    (cnu_pa_msg[202]),
	.first_din_203    (cnu_pa_msg[203]),
	.first_din_204    (cnu_pa_msg[204]),
	.first_din_205    (cnu_pa_msg[205]),
	.first_din_206    (cnu_pa_msg[206]),
	.first_din_207    (cnu_pa_msg[207]),
	.first_din_208    (cnu_pa_msg[208]),
	.first_din_209    (cnu_pa_msg[209]),
	.first_din_210    (cnu_pa_msg[210]),
	.first_din_211    (cnu_pa_msg[211]),
	.first_din_212    (cnu_pa_msg[212]),
	.first_din_213    (cnu_pa_msg[213]),
	.first_din_214    (cnu_pa_msg[214]),
	.first_din_215    (cnu_pa_msg[215]),
	.first_din_216    (cnu_pa_msg[216]),
	.first_din_217    (cnu_pa_msg[217]),
	.first_din_218    (cnu_pa_msg[218]),
	.first_din_219    (cnu_pa_msg[219]),
	.first_din_220    (cnu_pa_msg[220]),
	.first_din_221    (cnu_pa_msg[221]),
	.first_din_222    (cnu_pa_msg[222]),
	.first_din_223    (cnu_pa_msg[223]),
	.first_din_224    (cnu_pa_msg[224]),
	.first_din_225    (cnu_pa_msg[225]),
	.first_din_226    (cnu_pa_msg[226]),
	.first_din_227    (cnu_pa_msg[227]),
	.first_din_228    (cnu_pa_msg[228]),
	.first_din_229    (cnu_pa_msg[229]),
	.first_din_230    (cnu_pa_msg[230]),
	.first_din_231    (cnu_pa_msg[231]),
	.first_din_232    (cnu_pa_msg[232]),
	.first_din_233    (cnu_pa_msg[233]),
	.first_din_234    (cnu_pa_msg[234]),
	.first_din_235    (cnu_pa_msg[235]),
	.first_din_236    (cnu_pa_msg[236]),
	.first_din_237    (cnu_pa_msg[237]),
	.first_din_238    (cnu_pa_msg[238]),
	.first_din_239    (cnu_pa_msg[239]),
	.first_din_240    (cnu_pa_msg[240]),
	.first_din_241    (cnu_pa_msg[241]),
	.first_din_242    (cnu_pa_msg[242]),
	.first_din_243    (cnu_pa_msg[243]),
	.first_din_244    (cnu_pa_msg[244]),
	.first_din_245    (cnu_pa_msg[245]),
	.first_din_246    (cnu_pa_msg[246]),
	.first_din_247    (cnu_pa_msg[247]),
	.first_din_248    (cnu_pa_msg[248]),
	.first_din_249    (cnu_pa_msg[249]),
	.first_din_250    (cnu_pa_msg[250]),
	.first_din_251    (cnu_pa_msg[251]),
	.first_din_252    (cnu_pa_msg[252]),
	.first_din_253    (cnu_pa_msg[253]),
	.first_din_254    (cnu_pa_msg[254]),

	.second_din_0   (vnu_pa_msg[0]),
	.second_din_1   (vnu_pa_msg[1]),
	.second_din_2   (vnu_pa_msg[2]),
	.second_din_3   (vnu_pa_msg[3]),
	.second_din_4   (vnu_pa_msg[4]),
	.second_din_5   (vnu_pa_msg[5]),
	.second_din_6   (vnu_pa_msg[6]),
	.second_din_7   (vnu_pa_msg[7]),
	.second_din_8   (vnu_pa_msg[8]),
	.second_din_9   (vnu_pa_msg[9]),
	.second_din_10   (vnu_pa_msg[10]),
	.second_din_11   (vnu_pa_msg[11]),
	.second_din_12   (vnu_pa_msg[12]),
	.second_din_13   (vnu_pa_msg[13]),
	.second_din_14   (vnu_pa_msg[14]),
	.second_din_15   (vnu_pa_msg[15]),
	.second_din_16   (vnu_pa_msg[16]),
	.second_din_17   (vnu_pa_msg[17]),
	.second_din_18   (vnu_pa_msg[18]),
	.second_din_19   (vnu_pa_msg[19]),
	.second_din_20   (vnu_pa_msg[20]),
	.second_din_21   (vnu_pa_msg[21]),
	.second_din_22   (vnu_pa_msg[22]),
	.second_din_23   (vnu_pa_msg[23]),
	.second_din_24   (vnu_pa_msg[24]),
	.second_din_25   (vnu_pa_msg[25]),
	.second_din_26   (vnu_pa_msg[26]),
	.second_din_27   (vnu_pa_msg[27]),
	.second_din_28   (vnu_pa_msg[28]),
	.second_din_29   (vnu_pa_msg[29]),
	.second_din_30   (vnu_pa_msg[30]),
	.second_din_31   (vnu_pa_msg[31]),
	.second_din_32   (vnu_pa_msg[32]),
	.second_din_33   (vnu_pa_msg[33]),
	.second_din_34   (vnu_pa_msg[34]),
	.second_din_35   (vnu_pa_msg[35]),
	.second_din_36   (vnu_pa_msg[36]),
	.second_din_37   (vnu_pa_msg[37]),
	.second_din_38   (vnu_pa_msg[38]),
	.second_din_39   (vnu_pa_msg[39]),
	.second_din_40   (vnu_pa_msg[40]),
	.second_din_41   (vnu_pa_msg[41]),
	.second_din_42   (vnu_pa_msg[42]),
	.second_din_43   (vnu_pa_msg[43]),
	.second_din_44   (vnu_pa_msg[44]),
	.second_din_45   (vnu_pa_msg[45]),
	.second_din_46   (vnu_pa_msg[46]),
	.second_din_47   (vnu_pa_msg[47]),
	.second_din_48   (vnu_pa_msg[48]),
	.second_din_49   (vnu_pa_msg[49]),
	.second_din_50   (vnu_pa_msg[50]),
	.second_din_51   (vnu_pa_msg[51]),
	.second_din_52   (vnu_pa_msg[52]),
	.second_din_53   (vnu_pa_msg[53]),
	.second_din_54   (vnu_pa_msg[54]),
	.second_din_55   (vnu_pa_msg[55]),
	.second_din_56   (vnu_pa_msg[56]),
	.second_din_57   (vnu_pa_msg[57]),
	.second_din_58   (vnu_pa_msg[58]),
	.second_din_59   (vnu_pa_msg[59]),
	.second_din_60   (vnu_pa_msg[60]),
	.second_din_61   (vnu_pa_msg[61]),
	.second_din_62   (vnu_pa_msg[62]),
	.second_din_63   (vnu_pa_msg[63]),
	.second_din_64   (vnu_pa_msg[64]),
	.second_din_65   (vnu_pa_msg[65]),
	.second_din_66   (vnu_pa_msg[66]),
	.second_din_67   (vnu_pa_msg[67]),
	.second_din_68   (vnu_pa_msg[68]),
	.second_din_69   (vnu_pa_msg[69]),
	.second_din_70   (vnu_pa_msg[70]),
	.second_din_71   (vnu_pa_msg[71]),
	.second_din_72   (vnu_pa_msg[72]),
	.second_din_73   (vnu_pa_msg[73]),
	.second_din_74   (vnu_pa_msg[74]),
	.second_din_75   (vnu_pa_msg[75]),
	.second_din_76   (vnu_pa_msg[76]),
	.second_din_77   (vnu_pa_msg[77]),
	.second_din_78   (vnu_pa_msg[78]),
	.second_din_79   (vnu_pa_msg[79]),
	.second_din_80   (vnu_pa_msg[80]),
	.second_din_81   (vnu_pa_msg[81]),
	.second_din_82   (vnu_pa_msg[82]),
	.second_din_83   (vnu_pa_msg[83]),
	.second_din_84   (vnu_pa_msg[84]),
	.second_din_85   (vnu_pa_msg[85]),
	.second_din_86   (vnu_pa_msg[86]),
	.second_din_87   (vnu_pa_msg[87]),
	.second_din_88   (vnu_pa_msg[88]),
	.second_din_89   (vnu_pa_msg[89]),
	.second_din_90   (vnu_pa_msg[90]),
	.second_din_91   (vnu_pa_msg[91]),
	.second_din_92   (vnu_pa_msg[92]),
	.second_din_93   (vnu_pa_msg[93]),
	.second_din_94   (vnu_pa_msg[94]),
	.second_din_95   (vnu_pa_msg[95]),
	.second_din_96   (vnu_pa_msg[96]),
	.second_din_97   (vnu_pa_msg[97]),
	.second_din_98   (vnu_pa_msg[98]),
	.second_din_99   (vnu_pa_msg[99]),
	.second_din_100   (vnu_pa_msg[100]),
	.second_din_101   (vnu_pa_msg[101]),
	.second_din_102   (vnu_pa_msg[102]),
	.second_din_103   (vnu_pa_msg[103]),
	.second_din_104   (vnu_pa_msg[104]),
	.second_din_105   (vnu_pa_msg[105]),
	.second_din_106   (vnu_pa_msg[106]),
	.second_din_107   (vnu_pa_msg[107]),
	.second_din_108   (vnu_pa_msg[108]),
	.second_din_109   (vnu_pa_msg[109]),
	.second_din_110   (vnu_pa_msg[110]),
	.second_din_111   (vnu_pa_msg[111]),
	.second_din_112   (vnu_pa_msg[112]),
	.second_din_113   (vnu_pa_msg[113]),
	.second_din_114   (vnu_pa_msg[114]),
	.second_din_115   (vnu_pa_msg[115]),
	.second_din_116   (vnu_pa_msg[116]),
	.second_din_117   (vnu_pa_msg[117]),
	.second_din_118   (vnu_pa_msg[118]),
	.second_din_119   (vnu_pa_msg[119]),
	.second_din_120   (vnu_pa_msg[120]),
	.second_din_121   (vnu_pa_msg[121]),
	.second_din_122   (vnu_pa_msg[122]),
	.second_din_123   (vnu_pa_msg[123]),
	.second_din_124   (vnu_pa_msg[124]),
	.second_din_125   (vnu_pa_msg[125]),
	.second_din_126   (vnu_pa_msg[126]),
	.second_din_127   (vnu_pa_msg[127]),
	.second_din_128   (vnu_pa_msg[128]),
	.second_din_129   (vnu_pa_msg[129]),
	.second_din_130   (vnu_pa_msg[130]),
	.second_din_131   (vnu_pa_msg[131]),
	.second_din_132   (vnu_pa_msg[132]),
	.second_din_133   (vnu_pa_msg[133]),
	.second_din_134   (vnu_pa_msg[134]),
	.second_din_135   (vnu_pa_msg[135]),
	.second_din_136   (vnu_pa_msg[136]),
	.second_din_137   (vnu_pa_msg[137]),
	.second_din_138   (vnu_pa_msg[138]),
	.second_din_139   (vnu_pa_msg[139]),
	.second_din_140   (vnu_pa_msg[140]),
	.second_din_141   (vnu_pa_msg[141]),
	.second_din_142   (vnu_pa_msg[142]),
	.second_din_143   (vnu_pa_msg[143]),
	.second_din_144   (vnu_pa_msg[144]),
	.second_din_145   (vnu_pa_msg[145]),
	.second_din_146   (vnu_pa_msg[146]),
	.second_din_147   (vnu_pa_msg[147]),
	.second_din_148   (vnu_pa_msg[148]),
	.second_din_149   (vnu_pa_msg[149]),
	.second_din_150   (vnu_pa_msg[150]),
	.second_din_151   (vnu_pa_msg[151]),
	.second_din_152   (vnu_pa_msg[152]),
	.second_din_153   (vnu_pa_msg[153]),
	.second_din_154   (vnu_pa_msg[154]),
	.second_din_155   (vnu_pa_msg[155]),
	.second_din_156   (vnu_pa_msg[156]),
	.second_din_157   (vnu_pa_msg[157]),
	.second_din_158   (vnu_pa_msg[158]),
	.second_din_159   (vnu_pa_msg[159]),
	.second_din_160   (vnu_pa_msg[160]),
	.second_din_161   (vnu_pa_msg[161]),
	.second_din_162   (vnu_pa_msg[162]),
	.second_din_163   (vnu_pa_msg[163]),
	.second_din_164   (vnu_pa_msg[164]),
	.second_din_165   (vnu_pa_msg[165]),
	.second_din_166   (vnu_pa_msg[166]),
	.second_din_167   (vnu_pa_msg[167]),
	.second_din_168   (vnu_pa_msg[168]),
	.second_din_169   (vnu_pa_msg[169]),
	.second_din_170   (vnu_pa_msg[170]),
	.second_din_171   (vnu_pa_msg[171]),
	.second_din_172   (vnu_pa_msg[172]),
	.second_din_173   (vnu_pa_msg[173]),
	.second_din_174   (vnu_pa_msg[174]),
	.second_din_175   (vnu_pa_msg[175]),
	.second_din_176   (vnu_pa_msg[176]),
	.second_din_177   (vnu_pa_msg[177]),
	.second_din_178   (vnu_pa_msg[178]),
	.second_din_179   (vnu_pa_msg[179]),
	.second_din_180   (vnu_pa_msg[180]),
	.second_din_181   (vnu_pa_msg[181]),
	.second_din_182   (vnu_pa_msg[182]),
	.second_din_183   (vnu_pa_msg[183]),
	.second_din_184   (vnu_pa_msg[184]),
	.second_din_185   (vnu_pa_msg[185]),
	.second_din_186   (vnu_pa_msg[186]),
	.second_din_187   (vnu_pa_msg[187]),
	.second_din_188   (vnu_pa_msg[188]),
	.second_din_189   (vnu_pa_msg[189]),
	.second_din_190   (vnu_pa_msg[190]),
	.second_din_191   (vnu_pa_msg[191]),
	.second_din_192   (vnu_pa_msg[192]),
	.second_din_193   (vnu_pa_msg[193]),
	.second_din_194   (vnu_pa_msg[194]),
	.second_din_195   (vnu_pa_msg[195]),
	.second_din_196   (vnu_pa_msg[196]),
	.second_din_197   (vnu_pa_msg[197]),
	.second_din_198   (vnu_pa_msg[198]),
	.second_din_199   (vnu_pa_msg[199]),
	.second_din_200   (vnu_pa_msg[200]),
	.second_din_201   (vnu_pa_msg[201]),
	.second_din_202   (vnu_pa_msg[202]),
	.second_din_203   (vnu_pa_msg[203]),
	.second_din_204   (vnu_pa_msg[204]),
	.second_din_205   (vnu_pa_msg[205]),
	.second_din_206   (vnu_pa_msg[206]),
	.second_din_207   (vnu_pa_msg[207]),
	.second_din_208   (vnu_pa_msg[208]),
	.second_din_209   (vnu_pa_msg[209]),
	.second_din_210   (vnu_pa_msg[210]),
	.second_din_211   (vnu_pa_msg[211]),
	.second_din_212   (vnu_pa_msg[212]),
	.second_din_213   (vnu_pa_msg[213]),
	.second_din_214   (vnu_pa_msg[214]),
	.second_din_215   (vnu_pa_msg[215]),
	.second_din_216   (vnu_pa_msg[216]),
	.second_din_217   (vnu_pa_msg[217]),
	.second_din_218   (vnu_pa_msg[218]),
	.second_din_219   (vnu_pa_msg[219]),
	.second_din_220   (vnu_pa_msg[220]),
	.second_din_221   (vnu_pa_msg[221]),
	.second_din_222   (vnu_pa_msg[222]),
	.second_din_223   (vnu_pa_msg[223]),
	.second_din_224   (vnu_pa_msg[224]),
	.second_din_225   (vnu_pa_msg[225]),
	.second_din_226   (vnu_pa_msg[226]),
	.second_din_227   (vnu_pa_msg[227]),
	.second_din_228   (vnu_pa_msg[228]),
	.second_din_229   (vnu_pa_msg[229]),
	.second_din_230   (vnu_pa_msg[230]),
	.second_din_231   (vnu_pa_msg[231]),
	.second_din_232   (vnu_pa_msg[232]),
	.second_din_233   (vnu_pa_msg[233]),
	.second_din_234   (vnu_pa_msg[234]),
	.second_din_235   (vnu_pa_msg[235]),
	.second_din_236   (vnu_pa_msg[236]),
	.second_din_237   (vnu_pa_msg[237]),
	.second_din_238   (vnu_pa_msg[238]),
	.second_din_239   (vnu_pa_msg[239]),
	.second_din_240   (vnu_pa_msg[240]),
	.second_din_241   (vnu_pa_msg[241]),
	.second_din_242   (vnu_pa_msg[242]),
	.second_din_243   (vnu_pa_msg[243]),
	.second_din_244   (vnu_pa_msg[244]),
	.second_din_245   (vnu_pa_msg[245]),
	.second_din_246   (vnu_pa_msg[246]),
	.second_din_247   (vnu_pa_msg[247]),
	.second_din_248   (vnu_pa_msg[248]),
	.second_din_249   (vnu_pa_msg[249]),
	.second_din_250   (vnu_pa_msg[250]),
	.second_din_251   (vnu_pa_msg[251]),
	.second_din_252   (vnu_pa_msg[252]),
	.second_din_253   (vnu_pa_msg[253]),
	.second_din_254   (vnu_pa_msg[254]),

	.sync_addr_0    (cnu_sync_addr),
	.sync_addr_1    (vnu_sync_addr),
	.we             (we),
	.sys_clk        (sys_clk)
);
assign vnu_pa_msg_bit0[CHECK_PARALLELISM-1:0] = {vnu_pa_msg[254][0],vnu_pa_msg[253][0],vnu_pa_msg[252][0],vnu_pa_msg[251][0],vnu_pa_msg[250][0],vnu_pa_msg[249][0],vnu_pa_msg[248][0],vnu_pa_msg[247][0],vnu_pa_msg[246][0],vnu_pa_msg[245][0],vnu_pa_msg[244][0],vnu_pa_msg[243][0],vnu_pa_msg[242][0],vnu_pa_msg[241][0],vnu_pa_msg[240][0],vnu_pa_msg[239][0],vnu_pa_msg[238][0],vnu_pa_msg[237][0],vnu_pa_msg[236][0],vnu_pa_msg[235][0],vnu_pa_msg[234][0],vnu_pa_msg[233][0],vnu_pa_msg[232][0],vnu_pa_msg[231][0],vnu_pa_msg[230][0],vnu_pa_msg[229][0],vnu_pa_msg[228][0],vnu_pa_msg[227][0],vnu_pa_msg[226][0],vnu_pa_msg[225][0],vnu_pa_msg[224][0],vnu_pa_msg[223][0],vnu_pa_msg[222][0],vnu_pa_msg[221][0],vnu_pa_msg[220][0],vnu_pa_msg[219][0],vnu_pa_msg[218][0],vnu_pa_msg[217][0],vnu_pa_msg[216][0],vnu_pa_msg[215][0],vnu_pa_msg[214][0],vnu_pa_msg[213][0],vnu_pa_msg[212][0],vnu_pa_msg[211][0],vnu_pa_msg[210][0],vnu_pa_msg[209][0],vnu_pa_msg[208][0],vnu_pa_msg[207][0],vnu_pa_msg[206][0],vnu_pa_msg[205][0],vnu_pa_msg[204][0],vnu_pa_msg[203][0],vnu_pa_msg[202][0],vnu_pa_msg[201][0],vnu_pa_msg[200][0],vnu_pa_msg[199][0],vnu_pa_msg[198][0],vnu_pa_msg[197][0],vnu_pa_msg[196][0],vnu_pa_msg[195][0],vnu_pa_msg[194][0],vnu_pa_msg[193][0],vnu_pa_msg[192][0],vnu_pa_msg[191][0],vnu_pa_msg[190][0],vnu_pa_msg[189][0],vnu_pa_msg[188][0],vnu_pa_msg[187][0],vnu_pa_msg[186][0],vnu_pa_msg[185][0],vnu_pa_msg[184][0],vnu_pa_msg[183][0],vnu_pa_msg[182][0],vnu_pa_msg[181][0],vnu_pa_msg[180][0],vnu_pa_msg[179][0],vnu_pa_msg[178][0],vnu_pa_msg[177][0],vnu_pa_msg[176][0],vnu_pa_msg[175][0],vnu_pa_msg[174][0],vnu_pa_msg[173][0],vnu_pa_msg[172][0],vnu_pa_msg[171][0],vnu_pa_msg[170][0],vnu_pa_msg[169][0],vnu_pa_msg[168][0],vnu_pa_msg[167][0],vnu_pa_msg[166][0],vnu_pa_msg[165][0],vnu_pa_msg[164][0],vnu_pa_msg[163][0],vnu_pa_msg[162][0],vnu_pa_msg[161][0],vnu_pa_msg[160][0],vnu_pa_msg[159][0],vnu_pa_msg[158][0],vnu_pa_msg[157][0],vnu_pa_msg[156][0],vnu_pa_msg[155][0],vnu_pa_msg[154][0],vnu_pa_msg[153][0],vnu_pa_msg[152][0],vnu_pa_msg[151][0],vnu_pa_msg[150][0],vnu_pa_msg[149][0],vnu_pa_msg[148][0],vnu_pa_msg[147][0],vnu_pa_msg[146][0],vnu_pa_msg[145][0],vnu_pa_msg[144][0],vnu_pa_msg[143][0],vnu_pa_msg[142][0],vnu_pa_msg[141][0],vnu_pa_msg[140][0],vnu_pa_msg[139][0],vnu_pa_msg[138][0],vnu_pa_msg[137][0],vnu_pa_msg[136][0],vnu_pa_msg[135][0],vnu_pa_msg[134][0],vnu_pa_msg[133][0],vnu_pa_msg[132][0],vnu_pa_msg[131][0],vnu_pa_msg[130][0],vnu_pa_msg[129][0],vnu_pa_msg[128][0],vnu_pa_msg[127][0],vnu_pa_msg[126][0],vnu_pa_msg[125][0],vnu_pa_msg[124][0],vnu_pa_msg[123][0],vnu_pa_msg[122][0],vnu_pa_msg[121][0],vnu_pa_msg[120][0],vnu_pa_msg[119][0],vnu_pa_msg[118][0],vnu_pa_msg[117][0],vnu_pa_msg[116][0],vnu_pa_msg[115][0],vnu_pa_msg[114][0],vnu_pa_msg[113][0],vnu_pa_msg[112][0],vnu_pa_msg[111][0],vnu_pa_msg[110][0],vnu_pa_msg[109][0],vnu_pa_msg[108][0],vnu_pa_msg[107][0],vnu_pa_msg[106][0],vnu_pa_msg[105][0],vnu_pa_msg[104][0],vnu_pa_msg[103][0],vnu_pa_msg[102][0],vnu_pa_msg[101][0],vnu_pa_msg[100][0],vnu_pa_msg[99][0],vnu_pa_msg[98][0],vnu_pa_msg[97][0],vnu_pa_msg[96][0],vnu_pa_msg[95][0],vnu_pa_msg[94][0],vnu_pa_msg[93][0],vnu_pa_msg[92][0],vnu_pa_msg[91][0],vnu_pa_msg[90][0],vnu_pa_msg[89][0],vnu_pa_msg[88][0],vnu_pa_msg[87][0],vnu_pa_msg[86][0],vnu_pa_msg[85][0],vnu_pa_msg[84][0],vnu_pa_msg[83][0],vnu_pa_msg[82][0],vnu_pa_msg[81][0],vnu_pa_msg[80][0],vnu_pa_msg[79][0],vnu_pa_msg[78][0],vnu_pa_msg[77][0],vnu_pa_msg[76][0],vnu_pa_msg[75][0],vnu_pa_msg[74][0],vnu_pa_msg[73][0],vnu_pa_msg[72][0],vnu_pa_msg[71][0],vnu_pa_msg[70][0],vnu_pa_msg[69][0],vnu_pa_msg[68][0],vnu_pa_msg[67][0],vnu_pa_msg[66][0],vnu_pa_msg[65][0],vnu_pa_msg[64][0],vnu_pa_msg[63][0],vnu_pa_msg[62][0],vnu_pa_msg[61][0],vnu_pa_msg[60][0],vnu_pa_msg[59][0],vnu_pa_msg[58][0],vnu_pa_msg[57][0],vnu_pa_msg[56][0],vnu_pa_msg[55][0],vnu_pa_msg[54][0],vnu_pa_msg[53][0],vnu_pa_msg[52][0],vnu_pa_msg[51][0],vnu_pa_msg[50][0],vnu_pa_msg[49][0],vnu_pa_msg[48][0],vnu_pa_msg[47][0],vnu_pa_msg[46][0],vnu_pa_msg[45][0],vnu_pa_msg[44][0],vnu_pa_msg[43][0],vnu_pa_msg[42][0],vnu_pa_msg[41][0],vnu_pa_msg[40][0],vnu_pa_msg[39][0],vnu_pa_msg[38][0],vnu_pa_msg[37][0],vnu_pa_msg[36][0],vnu_pa_msg[35][0],vnu_pa_msg[34][0],vnu_pa_msg[33][0],vnu_pa_msg[32][0],vnu_pa_msg[31][0],vnu_pa_msg[30][0],vnu_pa_msg[29][0],vnu_pa_msg[28][0],vnu_pa_msg[27][0],vnu_pa_msg[26][0],vnu_pa_msg[25][0],vnu_pa_msg[24][0],vnu_pa_msg[23][0],vnu_pa_msg[22][0],vnu_pa_msg[21][0],vnu_pa_msg[20][0],vnu_pa_msg[19][0],vnu_pa_msg[18][0],vnu_pa_msg[17][0],vnu_pa_msg[16][0],vnu_pa_msg[15][0],vnu_pa_msg[14][0],vnu_pa_msg[13][0],vnu_pa_msg[12][0],vnu_pa_msg[11][0],vnu_pa_msg[10][0],vnu_pa_msg[9][0],vnu_pa_msg[8][0],vnu_pa_msg[7][0],vnu_pa_msg[6][0],vnu_pa_msg[5][0],vnu_pa_msg[4][0],vnu_pa_msg[3][0],vnu_pa_msg[2][0],vnu_pa_msg[1][0],vnu_pa_msg[0][0]};
assign pa_to_ch_ram[CH_DATA_WIDTH-1:0] = {vnu_pa_msg[254][QUAN_SIZE-1:0],vnu_pa_msg[253][QUAN_SIZE-1:0],vnu_pa_msg[252][QUAN_SIZE-1:0],vnu_pa_msg[251][QUAN_SIZE-1:0],vnu_pa_msg[250][QUAN_SIZE-1:0],vnu_pa_msg[249][QUAN_SIZE-1:0],vnu_pa_msg[248][QUAN_SIZE-1:0],vnu_pa_msg[247][QUAN_SIZE-1:0],vnu_pa_msg[246][QUAN_SIZE-1:0],vnu_pa_msg[245][QUAN_SIZE-1:0],vnu_pa_msg[244][QUAN_SIZE-1:0],vnu_pa_msg[243][QUAN_SIZE-1:0],vnu_pa_msg[242][QUAN_SIZE-1:0],vnu_pa_msg[241][QUAN_SIZE-1:0],vnu_pa_msg[240][QUAN_SIZE-1:0],vnu_pa_msg[239][QUAN_SIZE-1:0],vnu_pa_msg[238][QUAN_SIZE-1:0],vnu_pa_msg[237][QUAN_SIZE-1:0],vnu_pa_msg[236][QUAN_SIZE-1:0],vnu_pa_msg[235][QUAN_SIZE-1:0],vnu_pa_msg[234][QUAN_SIZE-1:0],vnu_pa_msg[233][QUAN_SIZE-1:0],vnu_pa_msg[232][QUAN_SIZE-1:0],vnu_pa_msg[231][QUAN_SIZE-1:0],vnu_pa_msg[230][QUAN_SIZE-1:0],vnu_pa_msg[229][QUAN_SIZE-1:0],vnu_pa_msg[228][QUAN_SIZE-1:0],vnu_pa_msg[227][QUAN_SIZE-1:0],vnu_pa_msg[226][QUAN_SIZE-1:0],vnu_pa_msg[225][QUAN_SIZE-1:0],vnu_pa_msg[224][QUAN_SIZE-1:0],vnu_pa_msg[223][QUAN_SIZE-1:0],vnu_pa_msg[222][QUAN_SIZE-1:0],vnu_pa_msg[221][QUAN_SIZE-1:0],vnu_pa_msg[220][QUAN_SIZE-1:0],vnu_pa_msg[219][QUAN_SIZE-1:0],vnu_pa_msg[218][QUAN_SIZE-1:0],vnu_pa_msg[217][QUAN_SIZE-1:0],vnu_pa_msg[216][QUAN_SIZE-1:0],vnu_pa_msg[215][QUAN_SIZE-1:0],vnu_pa_msg[214][QUAN_SIZE-1:0],vnu_pa_msg[213][QUAN_SIZE-1:0],vnu_pa_msg[212][QUAN_SIZE-1:0],vnu_pa_msg[211][QUAN_SIZE-1:0],vnu_pa_msg[210][QUAN_SIZE-1:0],vnu_pa_msg[209][QUAN_SIZE-1:0],vnu_pa_msg[208][QUAN_SIZE-1:0],vnu_pa_msg[207][QUAN_SIZE-1:0],vnu_pa_msg[206][QUAN_SIZE-1:0],vnu_pa_msg[205][QUAN_SIZE-1:0],vnu_pa_msg[204][QUAN_SIZE-1:0],vnu_pa_msg[203][QUAN_SIZE-1:0],vnu_pa_msg[202][QUAN_SIZE-1:0],vnu_pa_msg[201][QUAN_SIZE-1:0],vnu_pa_msg[200][QUAN_SIZE-1:0],vnu_pa_msg[199][QUAN_SIZE-1:0],vnu_pa_msg[198][QUAN_SIZE-1:0],vnu_pa_msg[197][QUAN_SIZE-1:0],vnu_pa_msg[196][QUAN_SIZE-1:0],vnu_pa_msg[195][QUAN_SIZE-1:0],vnu_pa_msg[194][QUAN_SIZE-1:0],vnu_pa_msg[193][QUAN_SIZE-1:0],vnu_pa_msg[192][QUAN_SIZE-1:0],vnu_pa_msg[191][QUAN_SIZE-1:0],vnu_pa_msg[190][QUAN_SIZE-1:0],vnu_pa_msg[189][QUAN_SIZE-1:0],vnu_pa_msg[188][QUAN_SIZE-1:0],vnu_pa_msg[187][QUAN_SIZE-1:0],vnu_pa_msg[186][QUAN_SIZE-1:0],vnu_pa_msg[185][QUAN_SIZE-1:0],vnu_pa_msg[184][QUAN_SIZE-1:0],vnu_pa_msg[183][QUAN_SIZE-1:0],vnu_pa_msg[182][QUAN_SIZE-1:0],vnu_pa_msg[181][QUAN_SIZE-1:0],vnu_pa_msg[180][QUAN_SIZE-1:0],vnu_pa_msg[179][QUAN_SIZE-1:0],vnu_pa_msg[178][QUAN_SIZE-1:0],vnu_pa_msg[177][QUAN_SIZE-1:0],vnu_pa_msg[176][QUAN_SIZE-1:0],vnu_pa_msg[175][QUAN_SIZE-1:0],vnu_pa_msg[174][QUAN_SIZE-1:0],vnu_pa_msg[173][QUAN_SIZE-1:0],vnu_pa_msg[172][QUAN_SIZE-1:0],vnu_pa_msg[171][QUAN_SIZE-1:0],vnu_pa_msg[170][QUAN_SIZE-1:0],vnu_pa_msg[169][QUAN_SIZE-1:0],vnu_pa_msg[168][QUAN_SIZE-1:0],vnu_pa_msg[167][QUAN_SIZE-1:0],vnu_pa_msg[166][QUAN_SIZE-1:0],vnu_pa_msg[165][QUAN_SIZE-1:0],vnu_pa_msg[164][QUAN_SIZE-1:0],vnu_pa_msg[163][QUAN_SIZE-1:0],vnu_pa_msg[162][QUAN_SIZE-1:0],vnu_pa_msg[161][QUAN_SIZE-1:0],vnu_pa_msg[160][QUAN_SIZE-1:0],vnu_pa_msg[159][QUAN_SIZE-1:0],vnu_pa_msg[158][QUAN_SIZE-1:0],vnu_pa_msg[157][QUAN_SIZE-1:0],vnu_pa_msg[156][QUAN_SIZE-1:0],vnu_pa_msg[155][QUAN_SIZE-1:0],vnu_pa_msg[154][QUAN_SIZE-1:0],vnu_pa_msg[153][QUAN_SIZE-1:0],vnu_pa_msg[152][QUAN_SIZE-1:0],vnu_pa_msg[151][QUAN_SIZE-1:0],vnu_pa_msg[150][QUAN_SIZE-1:0],vnu_pa_msg[149][QUAN_SIZE-1:0],vnu_pa_msg[148][QUAN_SIZE-1:0],vnu_pa_msg[147][QUAN_SIZE-1:0],vnu_pa_msg[146][QUAN_SIZE-1:0],vnu_pa_msg[145][QUAN_SIZE-1:0],vnu_pa_msg[144][QUAN_SIZE-1:0],vnu_pa_msg[143][QUAN_SIZE-1:0],vnu_pa_msg[142][QUAN_SIZE-1:0],vnu_pa_msg[141][QUAN_SIZE-1:0],vnu_pa_msg[140][QUAN_SIZE-1:0],vnu_pa_msg[139][QUAN_SIZE-1:0],vnu_pa_msg[138][QUAN_SIZE-1:0],vnu_pa_msg[137][QUAN_SIZE-1:0],vnu_pa_msg[136][QUAN_SIZE-1:0],vnu_pa_msg[135][QUAN_SIZE-1:0],vnu_pa_msg[134][QUAN_SIZE-1:0],vnu_pa_msg[133][QUAN_SIZE-1:0],vnu_pa_msg[132][QUAN_SIZE-1:0],vnu_pa_msg[131][QUAN_SIZE-1:0],vnu_pa_msg[130][QUAN_SIZE-1:0],vnu_pa_msg[129][QUAN_SIZE-1:0],vnu_pa_msg[128][QUAN_SIZE-1:0],vnu_pa_msg[127][QUAN_SIZE-1:0],vnu_pa_msg[126][QUAN_SIZE-1:0],vnu_pa_msg[125][QUAN_SIZE-1:0],vnu_pa_msg[124][QUAN_SIZE-1:0],vnu_pa_msg[123][QUAN_SIZE-1:0],vnu_pa_msg[122][QUAN_SIZE-1:0],vnu_pa_msg[121][QUAN_SIZE-1:0],vnu_pa_msg[120][QUAN_SIZE-1:0],vnu_pa_msg[119][QUAN_SIZE-1:0],vnu_pa_msg[118][QUAN_SIZE-1:0],vnu_pa_msg[117][QUAN_SIZE-1:0],vnu_pa_msg[116][QUAN_SIZE-1:0],vnu_pa_msg[115][QUAN_SIZE-1:0],vnu_pa_msg[114][QUAN_SIZE-1:0],vnu_pa_msg[113][QUAN_SIZE-1:0],vnu_pa_msg[112][QUAN_SIZE-1:0],vnu_pa_msg[111][QUAN_SIZE-1:0],vnu_pa_msg[110][QUAN_SIZE-1:0],vnu_pa_msg[109][QUAN_SIZE-1:0],vnu_pa_msg[108][QUAN_SIZE-1:0],vnu_pa_msg[107][QUAN_SIZE-1:0],vnu_pa_msg[106][QUAN_SIZE-1:0],vnu_pa_msg[105][QUAN_SIZE-1:0],vnu_pa_msg[104][QUAN_SIZE-1:0],vnu_pa_msg[103][QUAN_SIZE-1:0],vnu_pa_msg[102][QUAN_SIZE-1:0],vnu_pa_msg[101][QUAN_SIZE-1:0],vnu_pa_msg[100][QUAN_SIZE-1:0],vnu_pa_msg[99][QUAN_SIZE-1:0],vnu_pa_msg[98][QUAN_SIZE-1:0],vnu_pa_msg[97][QUAN_SIZE-1:0],vnu_pa_msg[96][QUAN_SIZE-1:0],vnu_pa_msg[95][QUAN_SIZE-1:0],vnu_pa_msg[94][QUAN_SIZE-1:0],vnu_pa_msg[93][QUAN_SIZE-1:0],vnu_pa_msg[92][QUAN_SIZE-1:0],vnu_pa_msg[91][QUAN_SIZE-1:0],vnu_pa_msg[90][QUAN_SIZE-1:0],vnu_pa_msg[89][QUAN_SIZE-1:0],vnu_pa_msg[88][QUAN_SIZE-1:0],vnu_pa_msg[87][QUAN_SIZE-1:0],vnu_pa_msg[86][QUAN_SIZE-1:0],vnu_pa_msg[85][QUAN_SIZE-1:0],vnu_pa_msg[84][QUAN_SIZE-1:0],vnu_pa_msg[83][QUAN_SIZE-1:0],vnu_pa_msg[82][QUAN_SIZE-1:0],vnu_pa_msg[81][QUAN_SIZE-1:0],vnu_pa_msg[80][QUAN_SIZE-1:0],vnu_pa_msg[79][QUAN_SIZE-1:0],vnu_pa_msg[78][QUAN_SIZE-1:0],vnu_pa_msg[77][QUAN_SIZE-1:0],vnu_pa_msg[76][QUAN_SIZE-1:0],vnu_pa_msg[75][QUAN_SIZE-1:0],vnu_pa_msg[74][QUAN_SIZE-1:0],vnu_pa_msg[73][QUAN_SIZE-1:0],vnu_pa_msg[72][QUAN_SIZE-1:0],vnu_pa_msg[71][QUAN_SIZE-1:0],vnu_pa_msg[70][QUAN_SIZE-1:0],vnu_pa_msg[69][QUAN_SIZE-1:0],vnu_pa_msg[68][QUAN_SIZE-1:0],vnu_pa_msg[67][QUAN_SIZE-1:0],vnu_pa_msg[66][QUAN_SIZE-1:0],vnu_pa_msg[65][QUAN_SIZE-1:0],vnu_pa_msg[64][QUAN_SIZE-1:0],vnu_pa_msg[63][QUAN_SIZE-1:0],vnu_pa_msg[62][QUAN_SIZE-1:0],vnu_pa_msg[61][QUAN_SIZE-1:0],vnu_pa_msg[60][QUAN_SIZE-1:0],vnu_pa_msg[59][QUAN_SIZE-1:0],vnu_pa_msg[58][QUAN_SIZE-1:0],vnu_pa_msg[57][QUAN_SIZE-1:0],vnu_pa_msg[56][QUAN_SIZE-1:0],vnu_pa_msg[55][QUAN_SIZE-1:0],vnu_pa_msg[54][QUAN_SIZE-1:0],vnu_pa_msg[53][QUAN_SIZE-1:0],vnu_pa_msg[52][QUAN_SIZE-1:0],vnu_pa_msg[51][QUAN_SIZE-1:0],vnu_pa_msg[50][QUAN_SIZE-1:0],vnu_pa_msg[49][QUAN_SIZE-1:0],vnu_pa_msg[48][QUAN_SIZE-1:0],vnu_pa_msg[47][QUAN_SIZE-1:0],vnu_pa_msg[46][QUAN_SIZE-1:0],vnu_pa_msg[45][QUAN_SIZE-1:0],vnu_pa_msg[44][QUAN_SIZE-1:0],vnu_pa_msg[43][QUAN_SIZE-1:0],vnu_pa_msg[42][QUAN_SIZE-1:0],vnu_pa_msg[41][QUAN_SIZE-1:0],vnu_pa_msg[40][QUAN_SIZE-1:0],vnu_pa_msg[39][QUAN_SIZE-1:0],vnu_pa_msg[38][QUAN_SIZE-1:0],vnu_pa_msg[37][QUAN_SIZE-1:0],vnu_pa_msg[36][QUAN_SIZE-1:0],vnu_pa_msg[35][QUAN_SIZE-1:0],vnu_pa_msg[34][QUAN_SIZE-1:0],vnu_pa_msg[33][QUAN_SIZE-1:0],vnu_pa_msg[32][QUAN_SIZE-1:0],vnu_pa_msg[31][QUAN_SIZE-1:0],vnu_pa_msg[30][QUAN_SIZE-1:0],vnu_pa_msg[29][QUAN_SIZE-1:0],vnu_pa_msg[28][QUAN_SIZE-1:0],vnu_pa_msg[27][QUAN_SIZE-1:0],vnu_pa_msg[26][QUAN_SIZE-1:0],vnu_pa_msg[25][QUAN_SIZE-1:0],vnu_pa_msg[24][QUAN_SIZE-1:0],vnu_pa_msg[23][QUAN_SIZE-1:0],vnu_pa_msg[22][QUAN_SIZE-1:0],vnu_pa_msg[21][QUAN_SIZE-1:0],vnu_pa_msg[20][QUAN_SIZE-1:0],vnu_pa_msg[19][QUAN_SIZE-1:0],vnu_pa_msg[18][QUAN_SIZE-1:0],vnu_pa_msg[17][QUAN_SIZE-1:0],vnu_pa_msg[16][QUAN_SIZE-1:0],vnu_pa_msg[15][QUAN_SIZE-1:0],vnu_pa_msg[14][QUAN_SIZE-1:0],vnu_pa_msg[13][QUAN_SIZE-1:0],vnu_pa_msg[12][QUAN_SIZE-1:0],vnu_pa_msg[11][QUAN_SIZE-1:0],vnu_pa_msg[10][QUAN_SIZE-1:0],vnu_pa_msg[9][QUAN_SIZE-1:0],vnu_pa_msg[8][QUAN_SIZE-1:0],vnu_pa_msg[7][QUAN_SIZE-1:0],vnu_pa_msg[6][QUAN_SIZE-1:0],vnu_pa_msg[5][QUAN_SIZE-1:0],vnu_pa_msg[4][QUAN_SIZE-1:0],vnu_pa_msg[3][QUAN_SIZE-1:0],vnu_pa_msg[2][QUAN_SIZE-1:0],vnu_pa_msg[1][QUAN_SIZE-1:0],vnu_pa_msg[0][QUAN_SIZE-1:0]};
endmodule
`endif