`include "define.vh"

`ifdef SCHED_4_6
module ram_pageAlign_interface_submatrix_7#(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 255,
	parameter LAYER_NUM = 3
) (
	output wire [QUAN_SIZE-1:0] msg_out_0,
	output wire [QUAN_SIZE-1:0] msg_out_1,
	output wire [QUAN_SIZE-1:0] msg_out_2,
	output wire [QUAN_SIZE-1:0] msg_out_3,
	output wire [QUAN_SIZE-1:0] msg_out_4,
	output wire [QUAN_SIZE-1:0] msg_out_5,
	output wire [QUAN_SIZE-1:0] msg_out_6,
	output wire [QUAN_SIZE-1:0] msg_out_7,
	output wire [QUAN_SIZE-1:0] msg_out_8,
	output wire [QUAN_SIZE-1:0] msg_out_9,
	output wire [QUAN_SIZE-1:0] msg_out_10,
	output wire [QUAN_SIZE-1:0] msg_out_11,
	output wire [QUAN_SIZE-1:0] msg_out_12,
	output wire [QUAN_SIZE-1:0] msg_out_13,
	output wire [QUAN_SIZE-1:0] msg_out_14,
	output wire [QUAN_SIZE-1:0] msg_out_15,
	output wire [QUAN_SIZE-1:0] msg_out_16,
	output wire [QUAN_SIZE-1:0] msg_out_17,
	output wire [QUAN_SIZE-1:0] msg_out_18,
	output wire [QUAN_SIZE-1:0] msg_out_19,
	output wire [QUAN_SIZE-1:0] msg_out_20,
	output wire [QUAN_SIZE-1:0] msg_out_21,
	output wire [QUAN_SIZE-1:0] msg_out_22,
	output wire [QUAN_SIZE-1:0] msg_out_23,
	output wire [QUAN_SIZE-1:0] msg_out_24,
	output wire [QUAN_SIZE-1:0] msg_out_25,
	output wire [QUAN_SIZE-1:0] msg_out_26,
	output wire [QUAN_SIZE-1:0] msg_out_27,
	output wire [QUAN_SIZE-1:0] msg_out_28,
	output wire [QUAN_SIZE-1:0] msg_out_29,
	output wire [QUAN_SIZE-1:0] msg_out_30,
	output wire [QUAN_SIZE-1:0] msg_out_31,
	output wire [QUAN_SIZE-1:0] msg_out_32,
	output wire [QUAN_SIZE-1:0] msg_out_33,
	output wire [QUAN_SIZE-1:0] msg_out_34,
	output wire [QUAN_SIZE-1:0] msg_out_35,
	output wire [QUAN_SIZE-1:0] msg_out_36,
	output wire [QUAN_SIZE-1:0] msg_out_37,
	output wire [QUAN_SIZE-1:0] msg_out_38,
	output wire [QUAN_SIZE-1:0] msg_out_39,
	output wire [QUAN_SIZE-1:0] msg_out_40,
	output wire [QUAN_SIZE-1:0] msg_out_41,
	output wire [QUAN_SIZE-1:0] msg_out_42,
	output wire [QUAN_SIZE-1:0] msg_out_43,
	output wire [QUAN_SIZE-1:0] msg_out_44,
	output wire [QUAN_SIZE-1:0] msg_out_45,
	output wire [QUAN_SIZE-1:0] msg_out_46,
	output wire [QUAN_SIZE-1:0] msg_out_47,
	output wire [QUAN_SIZE-1:0] msg_out_48,
	output wire [QUAN_SIZE-1:0] msg_out_49,
	output wire [QUAN_SIZE-1:0] msg_out_50,
	output wire [QUAN_SIZE-1:0] msg_out_51,
	output wire [QUAN_SIZE-1:0] msg_out_52,
	output wire [QUAN_SIZE-1:0] msg_out_53,
	output wire [QUAN_SIZE-1:0] msg_out_54,
	output wire [QUAN_SIZE-1:0] msg_out_55,
	output wire [QUAN_SIZE-1:0] msg_out_56,
	output wire [QUAN_SIZE-1:0] msg_out_57,
	output wire [QUAN_SIZE-1:0] msg_out_58,
	output wire [QUAN_SIZE-1:0] msg_out_59,
	output wire [QUAN_SIZE-1:0] msg_out_60,
	output wire [QUAN_SIZE-1:0] msg_out_61,
	output wire [QUAN_SIZE-1:0] msg_out_62,
	output wire [QUAN_SIZE-1:0] msg_out_63,
	output wire [QUAN_SIZE-1:0] msg_out_64,
	output wire [QUAN_SIZE-1:0] msg_out_65,
	output wire [QUAN_SIZE-1:0] msg_out_66,
	output wire [QUAN_SIZE-1:0] msg_out_67,
	output wire [QUAN_SIZE-1:0] msg_out_68,
	output wire [QUAN_SIZE-1:0] msg_out_69,
	output wire [QUAN_SIZE-1:0] msg_out_70,
	output wire [QUAN_SIZE-1:0] msg_out_71,
	output wire [QUAN_SIZE-1:0] msg_out_72,
	output wire [QUAN_SIZE-1:0] msg_out_73,
	output wire [QUAN_SIZE-1:0] msg_out_74,
	output wire [QUAN_SIZE-1:0] msg_out_75,
	output wire [QUAN_SIZE-1:0] msg_out_76,
	output wire [QUAN_SIZE-1:0] msg_out_77,
	output wire [QUAN_SIZE-1:0] msg_out_78,
	output wire [QUAN_SIZE-1:0] msg_out_79,
	output wire [QUAN_SIZE-1:0] msg_out_80,
	output wire [QUAN_SIZE-1:0] msg_out_81,
	output wire [QUAN_SIZE-1:0] msg_out_82,
	output wire [QUAN_SIZE-1:0] msg_out_83,
	output wire [QUAN_SIZE-1:0] msg_out_84,
	output wire [QUAN_SIZE-1:0] msg_out_85,
	output wire [QUAN_SIZE-1:0] msg_out_86,
	output wire [QUAN_SIZE-1:0] msg_out_87,
	output wire [QUAN_SIZE-1:0] msg_out_88,
	output wire [QUAN_SIZE-1:0] msg_out_89,
	output wire [QUAN_SIZE-1:0] msg_out_90,
	output wire [QUAN_SIZE-1:0] msg_out_91,
	output wire [QUAN_SIZE-1:0] msg_out_92,
	output wire [QUAN_SIZE-1:0] msg_out_93,
	output wire [QUAN_SIZE-1:0] msg_out_94,
	output wire [QUAN_SIZE-1:0] msg_out_95,
	output wire [QUAN_SIZE-1:0] msg_out_96,
	output wire [QUAN_SIZE-1:0] msg_out_97,
	output wire [QUAN_SIZE-1:0] msg_out_98,
	output wire [QUAN_SIZE-1:0] msg_out_99,
	output wire [QUAN_SIZE-1:0] msg_out_100,
	output wire [QUAN_SIZE-1:0] msg_out_101,
	output wire [QUAN_SIZE-1:0] msg_out_102,
	output wire [QUAN_SIZE-1:0] msg_out_103,
	output wire [QUAN_SIZE-1:0] msg_out_104,
	output wire [QUAN_SIZE-1:0] msg_out_105,
	output wire [QUAN_SIZE-1:0] msg_out_106,
	output wire [QUAN_SIZE-1:0] msg_out_107,
	output wire [QUAN_SIZE-1:0] msg_out_108,
	output wire [QUAN_SIZE-1:0] msg_out_109,
	output wire [QUAN_SIZE-1:0] msg_out_110,
	output wire [QUAN_SIZE-1:0] msg_out_111,
	output wire [QUAN_SIZE-1:0] msg_out_112,
	output wire [QUAN_SIZE-1:0] msg_out_113,
	output wire [QUAN_SIZE-1:0] msg_out_114,
	output wire [QUAN_SIZE-1:0] msg_out_115,
	output wire [QUAN_SIZE-1:0] msg_out_116,
	output wire [QUAN_SIZE-1:0] msg_out_117,
	output wire [QUAN_SIZE-1:0] msg_out_118,
	output wire [QUAN_SIZE-1:0] msg_out_119,
	output wire [QUAN_SIZE-1:0] msg_out_120,
	output wire [QUAN_SIZE-1:0] msg_out_121,
	output wire [QUAN_SIZE-1:0] msg_out_122,
	output wire [QUAN_SIZE-1:0] msg_out_123,
	output wire [QUAN_SIZE-1:0] msg_out_124,
	output wire [QUAN_SIZE-1:0] msg_out_125,
	output wire [QUAN_SIZE-1:0] msg_out_126,
	output wire [QUAN_SIZE-1:0] msg_out_127,
	output wire [QUAN_SIZE-1:0] msg_out_128,
	output wire [QUAN_SIZE-1:0] msg_out_129,
	output wire [QUAN_SIZE-1:0] msg_out_130,
	output wire [QUAN_SIZE-1:0] msg_out_131,
	output wire [QUAN_SIZE-1:0] msg_out_132,
	output wire [QUAN_SIZE-1:0] msg_out_133,
	output wire [QUAN_SIZE-1:0] msg_out_134,
	output wire [QUAN_SIZE-1:0] msg_out_135,
	output wire [QUAN_SIZE-1:0] msg_out_136,
	output wire [QUAN_SIZE-1:0] msg_out_137,
	output wire [QUAN_SIZE-1:0] msg_out_138,
	output wire [QUAN_SIZE-1:0] msg_out_139,
	output wire [QUAN_SIZE-1:0] msg_out_140,
	output wire [QUAN_SIZE-1:0] msg_out_141,
	output wire [QUAN_SIZE-1:0] msg_out_142,
	output wire [QUAN_SIZE-1:0] msg_out_143,
	output wire [QUAN_SIZE-1:0] msg_out_144,
	output wire [QUAN_SIZE-1:0] msg_out_145,
	output wire [QUAN_SIZE-1:0] msg_out_146,
	output wire [QUAN_SIZE-1:0] msg_out_147,
	output wire [QUAN_SIZE-1:0] msg_out_148,
	output wire [QUAN_SIZE-1:0] msg_out_149,
	output wire [QUAN_SIZE-1:0] msg_out_150,
	output wire [QUAN_SIZE-1:0] msg_out_151,
	output wire [QUAN_SIZE-1:0] msg_out_152,
	output wire [QUAN_SIZE-1:0] msg_out_153,
	output wire [QUAN_SIZE-1:0] msg_out_154,
	output wire [QUAN_SIZE-1:0] msg_out_155,
	output wire [QUAN_SIZE-1:0] msg_out_156,
	output wire [QUAN_SIZE-1:0] msg_out_157,
	output wire [QUAN_SIZE-1:0] msg_out_158,
	output wire [QUAN_SIZE-1:0] msg_out_159,
	output wire [QUAN_SIZE-1:0] msg_out_160,
	output wire [QUAN_SIZE-1:0] msg_out_161,
	output wire [QUAN_SIZE-1:0] msg_out_162,
	output wire [QUAN_SIZE-1:0] msg_out_163,
	output wire [QUAN_SIZE-1:0] msg_out_164,
	output wire [QUAN_SIZE-1:0] msg_out_165,
	output wire [QUAN_SIZE-1:0] msg_out_166,
	output wire [QUAN_SIZE-1:0] msg_out_167,
	output wire [QUAN_SIZE-1:0] msg_out_168,
	output wire [QUAN_SIZE-1:0] msg_out_169,
	output wire [QUAN_SIZE-1:0] msg_out_170,
	output wire [QUAN_SIZE-1:0] msg_out_171,
	output wire [QUAN_SIZE-1:0] msg_out_172,
	output wire [QUAN_SIZE-1:0] msg_out_173,
	output wire [QUAN_SIZE-1:0] msg_out_174,
	output wire [QUAN_SIZE-1:0] msg_out_175,
	output wire [QUAN_SIZE-1:0] msg_out_176,
	output wire [QUAN_SIZE-1:0] msg_out_177,
	output wire [QUAN_SIZE-1:0] msg_out_178,
	output wire [QUAN_SIZE-1:0] msg_out_179,
	output wire [QUAN_SIZE-1:0] msg_out_180,
	output wire [QUAN_SIZE-1:0] msg_out_181,
	output wire [QUAN_SIZE-1:0] msg_out_182,
	output wire [QUAN_SIZE-1:0] msg_out_183,
	output wire [QUAN_SIZE-1:0] msg_out_184,
	output wire [QUAN_SIZE-1:0] msg_out_185,
	output wire [QUAN_SIZE-1:0] msg_out_186,
	output wire [QUAN_SIZE-1:0] msg_out_187,
	output wire [QUAN_SIZE-1:0] msg_out_188,
	output wire [QUAN_SIZE-1:0] msg_out_189,
	output wire [QUAN_SIZE-1:0] msg_out_190,
	output wire [QUAN_SIZE-1:0] msg_out_191,
	output wire [QUAN_SIZE-1:0] msg_out_192,
	output wire [QUAN_SIZE-1:0] msg_out_193,
	output wire [QUAN_SIZE-1:0] msg_out_194,
	output wire [QUAN_SIZE-1:0] msg_out_195,
	output wire [QUAN_SIZE-1:0] msg_out_196,
	output wire [QUAN_SIZE-1:0] msg_out_197,
	output wire [QUAN_SIZE-1:0] msg_out_198,
	output wire [QUAN_SIZE-1:0] msg_out_199,
	output wire [QUAN_SIZE-1:0] msg_out_200,
	output wire [QUAN_SIZE-1:0] msg_out_201,
	output wire [QUAN_SIZE-1:0] msg_out_202,
	output wire [QUAN_SIZE-1:0] msg_out_203,
	output wire [QUAN_SIZE-1:0] msg_out_204,
	output wire [QUAN_SIZE-1:0] msg_out_205,
	output wire [QUAN_SIZE-1:0] msg_out_206,
	output wire [QUAN_SIZE-1:0] msg_out_207,
	output wire [QUAN_SIZE-1:0] msg_out_208,
	output wire [QUAN_SIZE-1:0] msg_out_209,
	output wire [QUAN_SIZE-1:0] msg_out_210,
	output wire [QUAN_SIZE-1:0] msg_out_211,
	output wire [QUAN_SIZE-1:0] msg_out_212,
	output wire [QUAN_SIZE-1:0] msg_out_213,
	output wire [QUAN_SIZE-1:0] msg_out_214,
	output wire [QUAN_SIZE-1:0] msg_out_215,
	output wire [QUAN_SIZE-1:0] msg_out_216,
	output wire [QUAN_SIZE-1:0] msg_out_217,
	output wire [QUAN_SIZE-1:0] msg_out_218,
	output wire [QUAN_SIZE-1:0] msg_out_219,
	output wire [QUAN_SIZE-1:0] msg_out_220,
	output wire [QUAN_SIZE-1:0] msg_out_221,
	output wire [QUAN_SIZE-1:0] msg_out_222,
	output wire [QUAN_SIZE-1:0] msg_out_223,
	output wire [QUAN_SIZE-1:0] msg_out_224,
	output wire [QUAN_SIZE-1:0] msg_out_225,
	output wire [QUAN_SIZE-1:0] msg_out_226,
	output wire [QUAN_SIZE-1:0] msg_out_227,
	output wire [QUAN_SIZE-1:0] msg_out_228,
	output wire [QUAN_SIZE-1:0] msg_out_229,
	output wire [QUAN_SIZE-1:0] msg_out_230,
	output wire [QUAN_SIZE-1:0] msg_out_231,
	output wire [QUAN_SIZE-1:0] msg_out_232,
	output wire [QUAN_SIZE-1:0] msg_out_233,
	output wire [QUAN_SIZE-1:0] msg_out_234,
	output wire [QUAN_SIZE-1:0] msg_out_235,
	output wire [QUAN_SIZE-1:0] msg_out_236,
	output wire [QUAN_SIZE-1:0] msg_out_237,
	output wire [QUAN_SIZE-1:0] msg_out_238,
	output wire [QUAN_SIZE-1:0] msg_out_239,
	output wire [QUAN_SIZE-1:0] msg_out_240,
	output wire [QUAN_SIZE-1:0] msg_out_241,
	output wire [QUAN_SIZE-1:0] msg_out_242,
	output wire [QUAN_SIZE-1:0] msg_out_243,
	output wire [QUAN_SIZE-1:0] msg_out_244,
	output wire [QUAN_SIZE-1:0] msg_out_245,
	output wire [QUAN_SIZE-1:0] msg_out_246,
	output wire [QUAN_SIZE-1:0] msg_out_247,
	output wire [QUAN_SIZE-1:0] msg_out_248,
	output wire [QUAN_SIZE-1:0] msg_out_249,
	output wire [QUAN_SIZE-1:0] msg_out_250,
	output wire [QUAN_SIZE-1:0] msg_out_251,
	output wire [QUAN_SIZE-1:0] msg_out_252,
	output wire [QUAN_SIZE-1:0] msg_out_253,
	output wire [QUAN_SIZE-1:0] msg_out_254,

	input wire [QUAN_SIZE-1:0] msg_in_0,
	input wire [QUAN_SIZE-1:0] msg_in_1,
	input wire [QUAN_SIZE-1:0] msg_in_2,
	input wire [QUAN_SIZE-1:0] msg_in_3,
	input wire [QUAN_SIZE-1:0] msg_in_4,
	input wire [QUAN_SIZE-1:0] msg_in_5,
	input wire [QUAN_SIZE-1:0] msg_in_6,
	input wire [QUAN_SIZE-1:0] msg_in_7,
	input wire [QUAN_SIZE-1:0] msg_in_8,
	input wire [QUAN_SIZE-1:0] msg_in_9,
	input wire [QUAN_SIZE-1:0] msg_in_10,
	input wire [QUAN_SIZE-1:0] msg_in_11,
	input wire [QUAN_SIZE-1:0] msg_in_12,
	input wire [QUAN_SIZE-1:0] msg_in_13,
	input wire [QUAN_SIZE-1:0] msg_in_14,
	input wire [QUAN_SIZE-1:0] msg_in_15,
	input wire [QUAN_SIZE-1:0] msg_in_16,
	input wire [QUAN_SIZE-1:0] msg_in_17,
	input wire [QUAN_SIZE-1:0] msg_in_18,
	input wire [QUAN_SIZE-1:0] msg_in_19,
	input wire [QUAN_SIZE-1:0] msg_in_20,
	input wire [QUAN_SIZE-1:0] msg_in_21,
	input wire [QUAN_SIZE-1:0] msg_in_22,
	input wire [QUAN_SIZE-1:0] msg_in_23,
	input wire [QUAN_SIZE-1:0] msg_in_24,
	input wire [QUAN_SIZE-1:0] msg_in_25,
	input wire [QUAN_SIZE-1:0] msg_in_26,
	input wire [QUAN_SIZE-1:0] msg_in_27,
	input wire [QUAN_SIZE-1:0] msg_in_28,
	input wire [QUAN_SIZE-1:0] msg_in_29,
	input wire [QUAN_SIZE-1:0] msg_in_30,
	input wire [QUAN_SIZE-1:0] msg_in_31,
	input wire [QUAN_SIZE-1:0] msg_in_32,
	input wire [QUAN_SIZE-1:0] msg_in_33,
	input wire [QUAN_SIZE-1:0] msg_in_34,
	input wire [QUAN_SIZE-1:0] msg_in_35,
	input wire [QUAN_SIZE-1:0] msg_in_36,
	input wire [QUAN_SIZE-1:0] msg_in_37,
	input wire [QUAN_SIZE-1:0] msg_in_38,
	input wire [QUAN_SIZE-1:0] msg_in_39,
	input wire [QUAN_SIZE-1:0] msg_in_40,
	input wire [QUAN_SIZE-1:0] msg_in_41,
	input wire [QUAN_SIZE-1:0] msg_in_42,
	input wire [QUAN_SIZE-1:0] msg_in_43,
	input wire [QUAN_SIZE-1:0] msg_in_44,
	input wire [QUAN_SIZE-1:0] msg_in_45,
	input wire [QUAN_SIZE-1:0] msg_in_46,
	input wire [QUAN_SIZE-1:0] msg_in_47,
	input wire [QUAN_SIZE-1:0] msg_in_48,
	input wire [QUAN_SIZE-1:0] msg_in_49,
	input wire [QUAN_SIZE-1:0] msg_in_50,
	input wire [QUAN_SIZE-1:0] msg_in_51,
	input wire [QUAN_SIZE-1:0] msg_in_52,
	input wire [QUAN_SIZE-1:0] msg_in_53,
	input wire [QUAN_SIZE-1:0] msg_in_54,
	input wire [QUAN_SIZE-1:0] msg_in_55,
	input wire [QUAN_SIZE-1:0] msg_in_56,
	input wire [QUAN_SIZE-1:0] msg_in_57,
	input wire [QUAN_SIZE-1:0] msg_in_58,
	input wire [QUAN_SIZE-1:0] msg_in_59,
	input wire [QUAN_SIZE-1:0] msg_in_60,
	input wire [QUAN_SIZE-1:0] msg_in_61,
	input wire [QUAN_SIZE-1:0] msg_in_62,
	input wire [QUAN_SIZE-1:0] msg_in_63,
	input wire [QUAN_SIZE-1:0] msg_in_64,
	input wire [QUAN_SIZE-1:0] msg_in_65,
	input wire [QUAN_SIZE-1:0] msg_in_66,
	input wire [QUAN_SIZE-1:0] msg_in_67,
	input wire [QUAN_SIZE-1:0] msg_in_68,
	input wire [QUAN_SIZE-1:0] msg_in_69,
	input wire [QUAN_SIZE-1:0] msg_in_70,
	input wire [QUAN_SIZE-1:0] msg_in_71,
	input wire [QUAN_SIZE-1:0] msg_in_72,
	input wire [QUAN_SIZE-1:0] msg_in_73,
	input wire [QUAN_SIZE-1:0] msg_in_74,
	input wire [QUAN_SIZE-1:0] msg_in_75,
	input wire [QUAN_SIZE-1:0] msg_in_76,
	input wire [QUAN_SIZE-1:0] msg_in_77,
	input wire [QUAN_SIZE-1:0] msg_in_78,
	input wire [QUAN_SIZE-1:0] msg_in_79,
	input wire [QUAN_SIZE-1:0] msg_in_80,
	input wire [QUAN_SIZE-1:0] msg_in_81,
	input wire [QUAN_SIZE-1:0] msg_in_82,
	input wire [QUAN_SIZE-1:0] msg_in_83,
	input wire [QUAN_SIZE-1:0] msg_in_84,
	input wire [QUAN_SIZE-1:0] msg_in_85,
	input wire [QUAN_SIZE-1:0] msg_in_86,
	input wire [QUAN_SIZE-1:0] msg_in_87,
	input wire [QUAN_SIZE-1:0] msg_in_88,
	input wire [QUAN_SIZE-1:0] msg_in_89,
	input wire [QUAN_SIZE-1:0] msg_in_90,
	input wire [QUAN_SIZE-1:0] msg_in_91,
	input wire [QUAN_SIZE-1:0] msg_in_92,
	input wire [QUAN_SIZE-1:0] msg_in_93,
	input wire [QUAN_SIZE-1:0] msg_in_94,
	input wire [QUAN_SIZE-1:0] msg_in_95,
	input wire [QUAN_SIZE-1:0] msg_in_96,
	input wire [QUAN_SIZE-1:0] msg_in_97,
	input wire [QUAN_SIZE-1:0] msg_in_98,
	input wire [QUAN_SIZE-1:0] msg_in_99,
	input wire [QUAN_SIZE-1:0] msg_in_100,
	input wire [QUAN_SIZE-1:0] msg_in_101,
	input wire [QUAN_SIZE-1:0] msg_in_102,
	input wire [QUAN_SIZE-1:0] msg_in_103,
	input wire [QUAN_SIZE-1:0] msg_in_104,
	input wire [QUAN_SIZE-1:0] msg_in_105,
	input wire [QUAN_SIZE-1:0] msg_in_106,
	input wire [QUAN_SIZE-1:0] msg_in_107,
	input wire [QUAN_SIZE-1:0] msg_in_108,
	input wire [QUAN_SIZE-1:0] msg_in_109,
	input wire [QUAN_SIZE-1:0] msg_in_110,
	input wire [QUAN_SIZE-1:0] msg_in_111,
	input wire [QUAN_SIZE-1:0] msg_in_112,
	input wire [QUAN_SIZE-1:0] msg_in_113,
	input wire [QUAN_SIZE-1:0] msg_in_114,
	input wire [QUAN_SIZE-1:0] msg_in_115,
	input wire [QUAN_SIZE-1:0] msg_in_116,
	input wire [QUAN_SIZE-1:0] msg_in_117,
	input wire [QUAN_SIZE-1:0] msg_in_118,
	input wire [QUAN_SIZE-1:0] msg_in_119,
	input wire [QUAN_SIZE-1:0] msg_in_120,
	input wire [QUAN_SIZE-1:0] msg_in_121,
	input wire [QUAN_SIZE-1:0] msg_in_122,
	input wire [QUAN_SIZE-1:0] msg_in_123,
	input wire [QUAN_SIZE-1:0] msg_in_124,
	input wire [QUAN_SIZE-1:0] msg_in_125,
	input wire [QUAN_SIZE-1:0] msg_in_126,
	input wire [QUAN_SIZE-1:0] msg_in_127,
	input wire [QUAN_SIZE-1:0] msg_in_128,
	input wire [QUAN_SIZE-1:0] msg_in_129,
	input wire [QUAN_SIZE-1:0] msg_in_130,
	input wire [QUAN_SIZE-1:0] msg_in_131,
	input wire [QUAN_SIZE-1:0] msg_in_132,
	input wire [QUAN_SIZE-1:0] msg_in_133,
	input wire [QUAN_SIZE-1:0] msg_in_134,
	input wire [QUAN_SIZE-1:0] msg_in_135,
	input wire [QUAN_SIZE-1:0] msg_in_136,
	input wire [QUAN_SIZE-1:0] msg_in_137,
	input wire [QUAN_SIZE-1:0] msg_in_138,
	input wire [QUAN_SIZE-1:0] msg_in_139,
	input wire [QUAN_SIZE-1:0] msg_in_140,
	input wire [QUAN_SIZE-1:0] msg_in_141,
	input wire [QUAN_SIZE-1:0] msg_in_142,
	input wire [QUAN_SIZE-1:0] msg_in_143,
	input wire [QUAN_SIZE-1:0] msg_in_144,
	input wire [QUAN_SIZE-1:0] msg_in_145,
	input wire [QUAN_SIZE-1:0] msg_in_146,
	input wire [QUAN_SIZE-1:0] msg_in_147,
	input wire [QUAN_SIZE-1:0] msg_in_148,
	input wire [QUAN_SIZE-1:0] msg_in_149,
	input wire [QUAN_SIZE-1:0] msg_in_150,
	input wire [QUAN_SIZE-1:0] msg_in_151,
	input wire [QUAN_SIZE-1:0] msg_in_152,
	input wire [QUAN_SIZE-1:0] msg_in_153,
	input wire [QUAN_SIZE-1:0] msg_in_154,
	input wire [QUAN_SIZE-1:0] msg_in_155,
	input wire [QUAN_SIZE-1:0] msg_in_156,
	input wire [QUAN_SIZE-1:0] msg_in_157,
	input wire [QUAN_SIZE-1:0] msg_in_158,
	input wire [QUAN_SIZE-1:0] msg_in_159,
	input wire [QUAN_SIZE-1:0] msg_in_160,
	input wire [QUAN_SIZE-1:0] msg_in_161,
	input wire [QUAN_SIZE-1:0] msg_in_162,
	input wire [QUAN_SIZE-1:0] msg_in_163,
	input wire [QUAN_SIZE-1:0] msg_in_164,
	input wire [QUAN_SIZE-1:0] msg_in_165,
	input wire [QUAN_SIZE-1:0] msg_in_166,
	input wire [QUAN_SIZE-1:0] msg_in_167,
	input wire [QUAN_SIZE-1:0] msg_in_168,
	input wire [QUAN_SIZE-1:0] msg_in_169,
	input wire [QUAN_SIZE-1:0] msg_in_170,
	input wire [QUAN_SIZE-1:0] msg_in_171,
	input wire [QUAN_SIZE-1:0] msg_in_172,
	input wire [QUAN_SIZE-1:0] msg_in_173,
	input wire [QUAN_SIZE-1:0] msg_in_174,
	input wire [QUAN_SIZE-1:0] msg_in_175,
	input wire [QUAN_SIZE-1:0] msg_in_176,
	input wire [QUAN_SIZE-1:0] msg_in_177,
	input wire [QUAN_SIZE-1:0] msg_in_178,
	input wire [QUAN_SIZE-1:0] msg_in_179,
	input wire [QUAN_SIZE-1:0] msg_in_180,
	input wire [QUAN_SIZE-1:0] msg_in_181,
	input wire [QUAN_SIZE-1:0] msg_in_182,
	input wire [QUAN_SIZE-1:0] msg_in_183,
	input wire [QUAN_SIZE-1:0] msg_in_184,
	input wire [QUAN_SIZE-1:0] msg_in_185,
	input wire [QUAN_SIZE-1:0] msg_in_186,
	input wire [QUAN_SIZE-1:0] msg_in_187,
	input wire [QUAN_SIZE-1:0] msg_in_188,
	input wire [QUAN_SIZE-1:0] msg_in_189,
	input wire [QUAN_SIZE-1:0] msg_in_190,
	input wire [QUAN_SIZE-1:0] msg_in_191,
	input wire [QUAN_SIZE-1:0] msg_in_192,
	input wire [QUAN_SIZE-1:0] msg_in_193,
	input wire [QUAN_SIZE-1:0] msg_in_194,
	input wire [QUAN_SIZE-1:0] msg_in_195,
	input wire [QUAN_SIZE-1:0] msg_in_196,
	input wire [QUAN_SIZE-1:0] msg_in_197,
	input wire [QUAN_SIZE-1:0] msg_in_198,
	input wire [QUAN_SIZE-1:0] msg_in_199,
	input wire [QUAN_SIZE-1:0] msg_in_200,
	input wire [QUAN_SIZE-1:0] msg_in_201,
	input wire [QUAN_SIZE-1:0] msg_in_202,
	input wire [QUAN_SIZE-1:0] msg_in_203,
	input wire [QUAN_SIZE-1:0] msg_in_204,
	input wire [QUAN_SIZE-1:0] msg_in_205,
	input wire [QUAN_SIZE-1:0] msg_in_206,
	input wire [QUAN_SIZE-1:0] msg_in_207,
	input wire [QUAN_SIZE-1:0] msg_in_208,
	input wire [QUAN_SIZE-1:0] msg_in_209,
	input wire [QUAN_SIZE-1:0] msg_in_210,
	input wire [QUAN_SIZE-1:0] msg_in_211,
	input wire [QUAN_SIZE-1:0] msg_in_212,
	input wire [QUAN_SIZE-1:0] msg_in_213,
	input wire [QUAN_SIZE-1:0] msg_in_214,
	input wire [QUAN_SIZE-1:0] msg_in_215,
	input wire [QUAN_SIZE-1:0] msg_in_216,
	input wire [QUAN_SIZE-1:0] msg_in_217,
	input wire [QUAN_SIZE-1:0] msg_in_218,
	input wire [QUAN_SIZE-1:0] msg_in_219,
	input wire [QUAN_SIZE-1:0] msg_in_220,
	input wire [QUAN_SIZE-1:0] msg_in_221,
	input wire [QUAN_SIZE-1:0] msg_in_222,
	input wire [QUAN_SIZE-1:0] msg_in_223,
	input wire [QUAN_SIZE-1:0] msg_in_224,
	input wire [QUAN_SIZE-1:0] msg_in_225,
	input wire [QUAN_SIZE-1:0] msg_in_226,
	input wire [QUAN_SIZE-1:0] msg_in_227,
	input wire [QUAN_SIZE-1:0] msg_in_228,
	input wire [QUAN_SIZE-1:0] msg_in_229,
	input wire [QUAN_SIZE-1:0] msg_in_230,
	input wire [QUAN_SIZE-1:0] msg_in_231,
	input wire [QUAN_SIZE-1:0] msg_in_232,
	input wire [QUAN_SIZE-1:0] msg_in_233,
	input wire [QUAN_SIZE-1:0] msg_in_234,
	input wire [QUAN_SIZE-1:0] msg_in_235,
	input wire [QUAN_SIZE-1:0] msg_in_236,
	input wire [QUAN_SIZE-1:0] msg_in_237,
	input wire [QUAN_SIZE-1:0] msg_in_238,
	input wire [QUAN_SIZE-1:0] msg_in_239,
	input wire [QUAN_SIZE-1:0] msg_in_240,
	input wire [QUAN_SIZE-1:0] msg_in_241,
	input wire [QUAN_SIZE-1:0] msg_in_242,
	input wire [QUAN_SIZE-1:0] msg_in_243,
	input wire [QUAN_SIZE-1:0] msg_in_244,
	input wire [QUAN_SIZE-1:0] msg_in_245,
	input wire [QUAN_SIZE-1:0] msg_in_246,
	input wire [QUAN_SIZE-1:0] msg_in_247,
	input wire [QUAN_SIZE-1:0] msg_in_248,
	input wire [QUAN_SIZE-1:0] msg_in_249,
	input wire [QUAN_SIZE-1:0] msg_in_250,
	input wire [QUAN_SIZE-1:0] msg_in_251,
	input wire [QUAN_SIZE-1:0] msg_in_252,
	input wire [QUAN_SIZE-1:0] msg_in_253,
	input wire [QUAN_SIZE-1:0] msg_in_254,

	input wire [LAYER_NUM-1:0] layer_status,
	input wire first_row_chunk,
	input wire sys_clk,
	input wire rstn
);

/////////////////////////////////////////////////////////////////////////////////////////////
// Main structure of Page Alignment Mechanism



/////////////////////////////////////////////////////////////////////////////////////////////
endmodule
`endif