`include "define.vh"

module fully_parallel_route(
	// (N-K) number of check-to-Variable message buses, each of which is d_c bit width as input ports of this routing network
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_00,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_01,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_02,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_03,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_04,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_05,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_10,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_11,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_12,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_13,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_14,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_15,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_20,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_21,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_22,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_23,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_24,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_25,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_30,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_31,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_32,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_33,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_34,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_35,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_40,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_41,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_42,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_43,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_44,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_45,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_50,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_51,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_52,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_53,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_54,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_55,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_60,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_61,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_62,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_63,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_64,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_65,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_70,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_71,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_72,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_73,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_74,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_75,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_80,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_81,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_82,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_83,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_84,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_85,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_90,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_91,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_92,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_93,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_94,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_95,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_100,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_101,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_102,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_103,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_104,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_105,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_110,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_111,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_112,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_113,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_114,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_115,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_120,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_121,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_122,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_123,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_124,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_125,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_130,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_131,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_132,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_133,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_134,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_135,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_140,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_141,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_142,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_143,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_144,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_145,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_150,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_151,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_152,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_153,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_154,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_155,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_160,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_161,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_162,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_163,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_164,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_165,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_170,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_171,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_172,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_173,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_174,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_175,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_180,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_181,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_182,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_183,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_184,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_185,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_190,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_191,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_192,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_193,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_194,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_195,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_200,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_201,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_202,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_203,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_204,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_205,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_210,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_211,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_212,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_213,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_214,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_215,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_220,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_221,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_222,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_223,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_224,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_225,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_230,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_231,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_232,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_233,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_234,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_235,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_240,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_241,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_242,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_243,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_244,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_245,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_250,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_251,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_252,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_253,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_254,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_255,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_260,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_261,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_262,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_263,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_264,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_265,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_270,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_271,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_272,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_273,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_274,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_275,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_280,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_281,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_282,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_283,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_284,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_285,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_290,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_291,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_292,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_293,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_294,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_295,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_300,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_301,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_302,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_303,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_304,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_305,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_310,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_311,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_312,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_313,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_314,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_315,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_320,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_321,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_322,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_323,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_324,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_325,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_330,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_331,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_332,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_333,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_334,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_335,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_340,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_341,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_342,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_343,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_344,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_345,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_350,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_351,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_352,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_353,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_354,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_355,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_360,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_361,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_362,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_363,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_364,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_365,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_370,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_371,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_372,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_373,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_374,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_375,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_380,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_381,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_382,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_383,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_384,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_385,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_390,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_391,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_392,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_393,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_394,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_395,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_400,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_401,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_402,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_403,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_404,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_405,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_410,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_411,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_412,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_413,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_414,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_415,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_420,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_421,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_422,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_423,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_424,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_425,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_430,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_431,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_432,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_433,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_434,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_435,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_440,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_441,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_442,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_443,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_444,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_445,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_450,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_451,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_452,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_453,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_454,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_455,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_460,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_461,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_462,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_463,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_464,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_465,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_470,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_471,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_472,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_473,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_474,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_475,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_480,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_481,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_482,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_483,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_484,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_485,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_490,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_491,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_492,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_493,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_494,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_495,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_500,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_501,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_502,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_503,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_504,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_505,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_510,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_511,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_512,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_513,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_514,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_515,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_520,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_521,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_522,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_523,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_524,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_525,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_530,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_531,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_532,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_533,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_534,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_535,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_540,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_541,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_542,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_543,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_544,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_545,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_550,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_551,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_552,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_553,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_554,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_555,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_560,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_561,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_562,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_563,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_564,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_565,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_570,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_571,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_572,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_573,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_574,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_575,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_580,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_581,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_582,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_583,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_584,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_585,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_590,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_591,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_592,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_593,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_594,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_595,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_600,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_601,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_602,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_603,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_604,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_605,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_610,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_611,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_612,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_613,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_614,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_615,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_620,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_621,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_622,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_623,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_624,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_625,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_630,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_631,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_632,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_633,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_634,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_635,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_640,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_641,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_642,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_643,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_644,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_645,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_650,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_651,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_652,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_653,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_654,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_655,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_660,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_661,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_662,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_663,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_664,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_665,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_670,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_671,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_672,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_673,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_674,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_675,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_680,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_681,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_682,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_683,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_684,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_685,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_690,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_691,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_692,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_693,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_694,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_695,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_700,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_701,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_702,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_703,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_704,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_705,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_710,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_711,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_712,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_713,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_714,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_715,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_720,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_721,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_722,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_723,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_724,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_725,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_730,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_731,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_732,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_733,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_734,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_735,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_740,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_741,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_742,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_743,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_744,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_745,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_750,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_751,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_752,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_753,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_754,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_755,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_760,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_761,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_762,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_763,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_764,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_765,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_770,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_771,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_772,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_773,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_774,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_775,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_780,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_781,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_782,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_783,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_784,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_785,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_790,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_791,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_792,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_793,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_794,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_795,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_800,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_801,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_802,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_803,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_804,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_805,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_810,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_811,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_812,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_813,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_814,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_815,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_820,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_821,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_822,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_823,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_824,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_825,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_830,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_831,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_832,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_833,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_834,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_835,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_840,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_841,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_842,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_843,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_844,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_845,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_850,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_851,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_852,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_853,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_854,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_855,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_860,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_861,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_862,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_863,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_864,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_865,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_870,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_871,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_872,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_873,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_874,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_875,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_880,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_881,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_882,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_883,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_884,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_885,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_890,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_891,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_892,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_893,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_894,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_895,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_900,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_901,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_902,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_903,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_904,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_905,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_910,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_911,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_912,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_913,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_914,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_915,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_920,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_921,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_922,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_923,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_924,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_925,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_930,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_931,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_932,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_933,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_934,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_935,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_940,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_941,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_942,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_943,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_944,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_945,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_950,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_951,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_952,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_953,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_954,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_955,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_960,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_961,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_962,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_963,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_964,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_965,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_970,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_971,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_972,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_973,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_974,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_975,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_980,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_981,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_982,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_983,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_984,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_985,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_990,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_991,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_992,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_993,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_994,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_995,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1000,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1001,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1002,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1003,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1004,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1005,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1010,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1011,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1012,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1013,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1014,
	output wire [`DATAPATH_WIDTH-1:0] v2c_parallelOut_1015,
	
	// N number of check-to-Variable message buses, each of which is d_v bit width outgoing to serial-to-parallel converters
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_00,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_01,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_02,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_10,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_11,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_12,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_20,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_21,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_22,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_30,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_31,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_32,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_40,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_41,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_42,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_50,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_51,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_52,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_60,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_61,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_62,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_70,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_71,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_72,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_80,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_81,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_82,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_90,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_91,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_92,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_100,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_101,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_102,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_110,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_111,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_112,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_120,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_121,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_122,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_130,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_131,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_132,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_140,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_141,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_142,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_150,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_151,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_152,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_160,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_161,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_162,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_170,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_171,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_172,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_180,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_181,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_182,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_190,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_191,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_192,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_200,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_201,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_202,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_210,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_211,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_212,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_220,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_221,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_222,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_230,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_231,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_232,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_240,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_241,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_242,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_250,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_251,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_252,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_260,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_261,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_262,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_270,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_271,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_272,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_280,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_281,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_282,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_290,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_291,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_292,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_300,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_301,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_302,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_310,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_311,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_312,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_320,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_321,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_322,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_330,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_331,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_332,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_340,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_341,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_342,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_350,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_351,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_352,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_360,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_361,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_362,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_370,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_371,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_372,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_380,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_381,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_382,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_390,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_391,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_392,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_400,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_401,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_402,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_410,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_411,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_412,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_420,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_421,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_422,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_430,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_431,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_432,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_440,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_441,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_442,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_450,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_451,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_452,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_460,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_461,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_462,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_470,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_471,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_472,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_480,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_481,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_482,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_490,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_491,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_492,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_500,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_501,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_502,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_510,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_511,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_512,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_520,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_521,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_522,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_530,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_531,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_532,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_540,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_541,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_542,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_550,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_551,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_552,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_560,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_561,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_562,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_570,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_571,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_572,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_580,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_581,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_582,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_590,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_591,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_592,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_600,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_601,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_602,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_610,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_611,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_612,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_620,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_621,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_622,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_630,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_631,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_632,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_640,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_641,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_642,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_650,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_651,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_652,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_660,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_661,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_662,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_670,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_671,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_672,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_680,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_681,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_682,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_690,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_691,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_692,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_700,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_701,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_702,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_710,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_711,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_712,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_720,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_721,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_722,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_730,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_731,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_732,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_740,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_741,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_742,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_750,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_751,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_752,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_760,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_761,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_762,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_770,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_771,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_772,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_780,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_781,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_782,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_790,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_791,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_792,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_800,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_801,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_802,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_810,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_811,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_812,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_820,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_821,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_822,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_830,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_831,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_832,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_840,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_841,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_842,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_850,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_851,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_852,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_860,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_861,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_862,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_870,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_871,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_872,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_880,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_881,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_882,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_890,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_891,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_892,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_900,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_901,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_902,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_910,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_911,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_912,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_920,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_921,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_922,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_930,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_931,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_932,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_940,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_941,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_942,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_950,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_951,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_952,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_960,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_961,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_962,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_970,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_971,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_972,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_980,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_981,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_982,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_990,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_991,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_992,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1000,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1001,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1002,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1010,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1011,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1012,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1020,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1021,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1022,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1030,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1031,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1032,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1040,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1041,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1042,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1050,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1051,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1052,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1060,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1061,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1062,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1070,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1071,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1072,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1080,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1081,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1082,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1090,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1091,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1092,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1100,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1101,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1102,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1110,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1111,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1112,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1120,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1121,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1122,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1130,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1131,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1132,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1140,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1141,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1142,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1150,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1151,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1152,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1160,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1161,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1162,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1170,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1171,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1172,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1180,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1181,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1182,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1190,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1191,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1192,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1200,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1201,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1202,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1210,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1211,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1212,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1220,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1221,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1222,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1230,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1231,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1232,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1240,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1241,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1242,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1250,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1251,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1252,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1260,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1261,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1262,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1270,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1271,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1272,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1280,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1281,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1282,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1290,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1291,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1292,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1300,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1301,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1302,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1310,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1311,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1312,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1320,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1321,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1322,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1330,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1331,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1332,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1340,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1341,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1342,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1350,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1351,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1352,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1360,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1361,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1362,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1370,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1371,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1372,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1380,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1381,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1382,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1390,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1391,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1392,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1400,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1401,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1402,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1410,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1411,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1412,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1420,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1421,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1422,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1430,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1431,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1432,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1440,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1441,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1442,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1450,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1451,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1452,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1460,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1461,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1462,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1470,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1471,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1472,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1480,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1481,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1482,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1490,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1491,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1492,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1500,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1501,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1502,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1510,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1511,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1512,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1520,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1521,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1522,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1530,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1531,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1532,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1540,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1541,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1542,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1550,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1551,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1552,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1560,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1561,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1562,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1570,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1571,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1572,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1580,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1581,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1582,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1590,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1591,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1592,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1600,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1601,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1602,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1610,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1611,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1612,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1620,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1621,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1622,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1630,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1631,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1632,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1640,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1641,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1642,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1650,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1651,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1652,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1660,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1661,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1662,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1670,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1671,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1672,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1680,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1681,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1682,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1690,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1691,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1692,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1700,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1701,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1702,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1710,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1711,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1712,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1720,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1721,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1722,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1730,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1731,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1732,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1740,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1741,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1742,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1750,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1751,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1752,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1760,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1761,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1762,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1770,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1771,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1772,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1780,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1781,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1782,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1790,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1791,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1792,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1800,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1801,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1802,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1810,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1811,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1812,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1820,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1821,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1822,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1830,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1831,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1832,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1840,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1841,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1842,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1850,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1851,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1852,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1860,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1861,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1862,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1870,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1871,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1872,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1880,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1881,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1882,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1890,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1891,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1892,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1900,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1901,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1902,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1910,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1911,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1912,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1920,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1921,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1922,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1930,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1931,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1932,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1940,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1941,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1942,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1950,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1951,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1952,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1960,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1961,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1962,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1970,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1971,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1972,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1980,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1981,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1982,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1990,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1991,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_1992,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2000,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2001,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2002,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2010,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2011,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2012,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2020,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2021,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2022,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2030,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2031,
	output wire [`DATAPATH_WIDTH-1:0] c2v_parallelOut_2032,
	
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_00,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_01,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_02,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_03,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_04,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_05,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_10,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_11,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_12,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_13,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_14,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_15,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_20,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_21,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_22,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_23,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_24,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_25,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_30,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_31,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_32,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_33,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_34,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_35,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_40,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_41,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_42,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_43,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_44,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_45,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_50,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_51,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_52,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_53,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_54,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_55,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_60,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_61,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_62,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_63,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_64,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_65,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_70,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_71,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_72,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_73,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_74,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_75,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_80,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_81,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_82,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_83,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_84,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_85,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_90,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_91,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_92,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_93,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_94,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_95,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_100,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_101,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_102,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_103,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_104,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_105,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_110,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_111,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_112,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_113,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_114,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_115,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_120,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_121,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_122,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_123,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_124,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_125,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_130,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_131,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_132,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_133,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_134,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_135,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_140,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_141,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_142,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_143,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_144,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_145,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_150,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_151,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_152,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_153,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_154,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_155,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_160,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_161,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_162,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_163,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_164,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_165,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_170,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_171,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_172,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_173,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_174,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_175,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_180,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_181,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_182,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_183,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_184,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_185,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_190,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_191,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_192,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_193,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_194,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_195,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_200,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_201,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_202,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_203,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_204,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_205,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_210,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_211,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_212,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_213,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_214,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_215,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_220,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_221,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_222,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_223,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_224,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_225,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_230,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_231,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_232,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_233,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_234,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_235,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_240,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_241,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_242,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_243,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_244,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_245,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_250,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_251,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_252,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_253,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_254,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_255,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_260,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_261,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_262,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_263,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_264,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_265,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_270,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_271,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_272,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_273,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_274,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_275,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_280,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_281,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_282,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_283,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_284,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_285,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_290,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_291,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_292,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_293,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_294,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_295,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_300,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_301,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_302,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_303,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_304,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_305,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_310,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_311,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_312,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_313,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_314,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_315,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_320,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_321,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_322,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_323,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_324,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_325,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_330,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_331,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_332,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_333,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_334,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_335,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_340,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_341,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_342,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_343,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_344,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_345,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_350,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_351,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_352,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_353,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_354,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_355,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_360,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_361,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_362,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_363,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_364,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_365,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_370,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_371,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_372,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_373,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_374,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_375,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_380,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_381,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_382,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_383,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_384,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_385,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_390,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_391,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_392,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_393,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_394,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_395,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_400,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_401,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_402,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_403,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_404,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_405,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_410,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_411,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_412,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_413,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_414,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_415,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_420,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_421,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_422,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_423,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_424,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_425,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_430,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_431,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_432,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_433,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_434,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_435,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_440,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_441,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_442,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_443,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_444,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_445,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_450,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_451,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_452,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_453,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_454,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_455,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_460,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_461,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_462,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_463,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_464,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_465,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_470,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_471,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_472,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_473,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_474,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_475,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_480,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_481,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_482,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_483,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_484,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_485,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_490,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_491,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_492,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_493,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_494,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_495,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_500,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_501,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_502,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_503,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_504,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_505,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_510,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_511,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_512,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_513,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_514,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_515,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_520,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_521,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_522,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_523,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_524,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_525,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_530,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_531,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_532,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_533,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_534,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_535,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_540,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_541,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_542,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_543,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_544,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_545,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_550,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_551,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_552,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_553,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_554,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_555,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_560,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_561,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_562,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_563,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_564,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_565,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_570,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_571,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_572,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_573,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_574,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_575,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_580,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_581,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_582,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_583,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_584,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_585,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_590,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_591,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_592,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_593,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_594,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_595,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_600,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_601,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_602,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_603,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_604,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_605,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_610,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_611,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_612,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_613,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_614,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_615,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_620,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_621,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_622,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_623,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_624,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_625,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_630,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_631,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_632,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_633,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_634,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_635,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_640,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_641,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_642,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_643,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_644,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_645,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_650,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_651,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_652,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_653,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_654,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_655,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_660,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_661,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_662,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_663,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_664,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_665,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_670,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_671,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_672,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_673,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_674,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_675,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_680,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_681,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_682,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_683,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_684,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_685,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_690,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_691,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_692,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_693,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_694,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_695,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_700,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_701,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_702,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_703,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_704,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_705,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_710,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_711,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_712,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_713,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_714,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_715,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_720,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_721,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_722,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_723,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_724,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_725,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_730,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_731,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_732,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_733,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_734,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_735,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_740,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_741,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_742,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_743,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_744,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_745,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_750,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_751,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_752,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_753,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_754,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_755,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_760,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_761,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_762,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_763,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_764,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_765,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_770,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_771,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_772,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_773,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_774,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_775,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_780,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_781,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_782,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_783,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_784,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_785,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_790,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_791,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_792,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_793,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_794,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_795,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_800,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_801,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_802,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_803,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_804,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_805,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_810,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_811,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_812,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_813,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_814,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_815,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_820,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_821,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_822,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_823,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_824,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_825,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_830,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_831,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_832,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_833,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_834,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_835,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_840,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_841,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_842,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_843,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_844,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_845,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_850,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_851,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_852,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_853,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_854,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_855,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_860,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_861,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_862,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_863,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_864,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_865,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_870,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_871,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_872,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_873,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_874,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_875,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_880,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_881,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_882,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_883,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_884,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_885,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_890,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_891,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_892,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_893,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_894,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_895,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_900,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_901,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_902,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_903,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_904,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_905,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_910,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_911,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_912,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_913,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_914,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_915,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_920,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_921,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_922,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_923,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_924,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_925,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_930,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_931,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_932,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_933,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_934,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_935,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_940,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_941,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_942,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_943,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_944,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_945,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_950,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_951,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_952,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_953,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_954,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_955,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_960,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_961,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_962,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_963,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_964,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_965,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_970,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_971,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_972,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_973,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_974,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_975,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_980,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_981,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_982,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_983,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_984,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_985,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_990,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_991,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_992,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_993,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_994,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_995,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1000,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1001,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1002,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1003,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1004,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1005,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1010,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1011,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1012,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1013,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1014,
	input wire [`DATAPATH_WIDTH-1:0] c2v_parallelIn_1015,
	
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_00,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_01,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_02,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_10,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_11,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_12,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_20,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_21,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_22,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_30,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_31,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_32,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_40,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_41,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_42,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_50,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_51,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_52,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_60,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_61,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_62,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_70,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_71,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_72,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_80,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_81,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_82,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_90,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_91,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_92,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_100,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_101,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_102,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_110,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_111,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_112,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_120,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_121,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_122,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_130,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_131,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_132,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_140,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_141,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_142,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_150,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_151,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_152,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_160,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_161,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_162,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_170,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_171,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_172,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_180,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_181,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_182,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_190,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_191,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_192,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_200,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_201,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_202,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_210,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_211,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_212,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_220,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_221,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_222,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_230,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_231,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_232,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_240,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_241,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_242,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_250,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_251,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_252,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_260,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_261,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_262,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_270,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_271,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_272,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_280,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_281,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_282,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_290,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_291,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_292,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_300,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_301,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_302,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_310,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_311,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_312,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_320,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_321,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_322,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_330,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_331,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_332,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_340,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_341,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_342,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_350,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_351,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_352,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_360,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_361,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_362,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_370,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_371,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_372,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_380,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_381,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_382,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_390,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_391,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_392,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_400,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_401,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_402,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_410,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_411,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_412,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_420,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_421,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_422,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_430,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_431,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_432,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_440,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_441,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_442,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_450,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_451,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_452,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_460,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_461,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_462,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_470,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_471,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_472,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_480,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_481,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_482,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_490,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_491,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_492,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_500,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_501,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_502,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_510,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_511,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_512,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_520,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_521,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_522,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_530,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_531,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_532,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_540,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_541,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_542,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_550,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_551,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_552,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_560,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_561,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_562,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_570,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_571,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_572,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_580,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_581,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_582,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_590,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_591,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_592,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_600,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_601,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_602,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_610,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_611,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_612,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_620,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_621,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_622,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_630,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_631,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_632,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_640,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_641,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_642,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_650,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_651,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_652,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_660,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_661,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_662,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_670,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_671,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_672,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_680,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_681,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_682,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_690,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_691,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_692,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_700,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_701,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_702,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_710,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_711,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_712,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_720,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_721,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_722,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_730,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_731,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_732,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_740,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_741,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_742,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_750,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_751,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_752,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_760,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_761,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_762,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_770,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_771,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_772,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_780,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_781,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_782,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_790,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_791,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_792,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_800,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_801,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_802,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_810,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_811,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_812,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_820,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_821,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_822,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_830,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_831,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_832,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_840,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_841,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_842,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_850,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_851,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_852,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_860,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_861,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_862,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_870,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_871,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_872,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_880,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_881,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_882,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_890,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_891,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_892,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_900,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_901,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_902,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_910,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_911,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_912,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_920,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_921,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_922,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_930,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_931,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_932,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_940,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_941,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_942,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_950,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_951,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_952,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_960,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_961,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_962,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_970,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_971,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_972,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_980,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_981,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_982,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_990,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_991,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_992,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1000,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1001,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1002,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1010,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1011,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1012,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1020,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1021,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1022,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1030,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1031,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1032,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1040,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1041,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1042,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1050,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1051,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1052,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1060,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1061,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1062,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1070,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1071,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1072,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1080,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1081,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1082,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1090,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1091,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1092,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1100,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1101,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1102,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1110,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1111,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1112,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1120,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1121,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1122,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1130,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1131,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1132,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1140,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1141,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1142,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1150,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1151,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1152,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1160,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1161,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1162,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1170,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1171,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1172,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1180,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1181,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1182,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1190,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1191,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1192,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1200,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1201,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1202,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1210,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1211,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1212,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1220,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1221,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1222,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1230,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1231,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1232,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1240,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1241,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1242,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1250,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1251,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1252,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1260,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1261,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1262,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1270,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1271,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1272,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1280,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1281,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1282,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1290,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1291,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1292,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1300,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1301,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1302,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1310,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1311,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1312,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1320,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1321,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1322,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1330,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1331,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1332,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1340,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1341,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1342,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1350,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1351,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1352,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1360,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1361,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1362,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1370,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1371,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1372,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1380,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1381,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1382,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1390,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1391,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1392,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1400,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1401,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1402,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1410,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1411,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1412,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1420,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1421,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1422,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1430,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1431,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1432,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1440,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1441,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1442,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1450,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1451,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1452,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1460,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1461,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1462,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1470,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1471,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1472,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1480,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1481,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1482,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1490,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1491,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1492,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1500,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1501,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1502,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1510,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1511,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1512,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1520,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1521,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1522,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1530,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1531,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1532,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1540,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1541,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1542,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1550,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1551,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1552,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1560,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1561,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1562,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1570,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1571,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1572,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1580,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1581,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1582,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1590,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1591,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1592,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1600,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1601,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1602,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1610,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1611,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1612,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1620,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1621,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1622,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1630,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1631,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1632,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1640,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1641,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1642,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1650,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1651,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1652,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1660,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1661,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1662,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1670,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1671,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1672,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1680,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1681,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1682,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1690,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1691,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1692,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1700,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1701,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1702,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1710,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1711,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1712,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1720,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1721,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1722,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1730,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1731,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1732,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1740,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1741,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1742,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1750,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1751,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1752,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1760,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1761,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1762,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1770,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1771,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1772,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1780,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1781,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1782,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1790,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1791,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1792,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1800,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1801,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1802,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1810,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1811,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1812,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1820,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1821,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1822,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1830,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1831,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1832,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1840,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1841,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1842,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1850,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1851,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1852,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1860,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1861,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1862,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1870,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1871,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1872,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1880,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1881,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1882,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1890,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1891,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1892,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1900,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1901,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1902,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1910,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1911,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1912,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1920,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1921,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1922,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1930,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1931,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1932,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1940,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1941,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1942,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1950,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1951,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1952,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1960,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1961,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1962,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1970,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1971,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1972,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1980,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1981,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1982,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1990,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1991,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_1992,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2000,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2001,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2002,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2010,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2011,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2012,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2020,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2021,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2022,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2030,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2031,
	input wire [`DATAPATH_WIDTH-1:0] v2c_parallelIn_2032,
	
	input wire [1:0] load,
	input wire [1:0] parallel_en,
	input wire serial_clk
);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_0;
	cnu_bitSerial_port cnu_converter_port0(
		.serialInOut (cn_serialInOut_0[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_00[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_01[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_02[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_03[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_04[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_05[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_00[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_01[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_02[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_03[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_04[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_05[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_1;
	cnu_bitSerial_port cnu_converter_port1(
		.serialInOut (cn_serialInOut_1[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_10[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_11[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_12[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_13[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_14[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_15[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_10[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_11[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_12[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_13[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_14[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_15[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_2;
	cnu_bitSerial_port cnu_converter_port2(
		.serialInOut (cn_serialInOut_2[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_20[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_21[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_22[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_23[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_24[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_25[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_20[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_21[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_22[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_23[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_24[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_25[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_3;
	cnu_bitSerial_port cnu_converter_port3(
		.serialInOut (cn_serialInOut_3[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_30[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_31[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_32[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_33[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_34[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_35[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_30[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_31[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_32[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_33[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_34[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_35[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_4;
	cnu_bitSerial_port cnu_converter_port4(
		.serialInOut (cn_serialInOut_4[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_40[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_41[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_42[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_43[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_44[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_45[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_40[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_41[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_42[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_43[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_44[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_45[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_5;
	cnu_bitSerial_port cnu_converter_port5(
		.serialInOut (cn_serialInOut_5[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_50[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_51[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_52[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_53[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_54[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_55[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_50[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_51[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_52[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_53[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_54[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_55[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_6;
	cnu_bitSerial_port cnu_converter_port6(
		.serialInOut (cn_serialInOut_6[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_60[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_61[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_62[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_63[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_64[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_65[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_60[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_61[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_62[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_63[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_64[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_65[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_7;
	cnu_bitSerial_port cnu_converter_port7(
		.serialInOut (cn_serialInOut_7[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_70[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_71[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_72[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_73[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_74[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_75[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_70[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_71[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_72[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_73[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_74[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_75[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_8;
	cnu_bitSerial_port cnu_converter_port8(
		.serialInOut (cn_serialInOut_8[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_80[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_81[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_82[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_83[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_84[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_85[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_80[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_81[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_82[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_83[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_84[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_85[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_9;
	cnu_bitSerial_port cnu_converter_port9(
		.serialInOut (cn_serialInOut_9[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_90[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_91[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_92[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_93[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_94[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_95[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_90[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_91[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_92[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_93[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_94[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_95[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_10;
	cnu_bitSerial_port cnu_converter_port10(
		.serialInOut (cn_serialInOut_10[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_100[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_101[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_102[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_103[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_104[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_105[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_100[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_101[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_102[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_103[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_104[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_105[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_11;
	cnu_bitSerial_port cnu_converter_port11(
		.serialInOut (cn_serialInOut_11[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_110[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_111[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_112[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_113[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_114[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_115[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_110[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_111[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_112[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_113[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_114[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_115[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_12;
	cnu_bitSerial_port cnu_converter_port12(
		.serialInOut (cn_serialInOut_12[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_120[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_121[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_122[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_123[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_124[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_125[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_120[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_121[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_122[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_123[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_124[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_125[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_13;
	cnu_bitSerial_port cnu_converter_port13(
		.serialInOut (cn_serialInOut_13[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_130[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_131[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_132[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_133[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_134[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_135[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_130[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_131[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_132[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_133[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_134[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_135[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_14;
	cnu_bitSerial_port cnu_converter_port14(
		.serialInOut (cn_serialInOut_14[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_140[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_141[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_142[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_143[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_144[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_145[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_140[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_141[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_142[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_143[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_144[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_145[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_15;
	cnu_bitSerial_port cnu_converter_port15(
		.serialInOut (cn_serialInOut_15[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_150[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_151[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_152[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_153[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_154[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_155[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_150[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_151[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_152[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_153[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_154[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_155[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_16;
	cnu_bitSerial_port cnu_converter_port16(
		.serialInOut (cn_serialInOut_16[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_160[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_161[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_162[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_163[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_164[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_165[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_160[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_161[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_162[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_163[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_164[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_165[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_17;
	cnu_bitSerial_port cnu_converter_port17(
		.serialInOut (cn_serialInOut_17[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_170[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_171[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_172[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_173[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_174[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_175[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_170[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_171[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_172[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_173[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_174[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_175[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_18;
	cnu_bitSerial_port cnu_converter_port18(
		.serialInOut (cn_serialInOut_18[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_180[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_181[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_182[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_183[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_184[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_185[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_180[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_181[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_182[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_183[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_184[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_185[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_19;
	cnu_bitSerial_port cnu_converter_port19(
		.serialInOut (cn_serialInOut_19[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_190[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_191[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_192[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_193[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_194[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_195[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_190[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_191[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_192[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_193[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_194[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_195[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_20;
	cnu_bitSerial_port cnu_converter_port20(
		.serialInOut (cn_serialInOut_20[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_200[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_201[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_202[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_203[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_204[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_205[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_200[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_201[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_202[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_203[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_204[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_205[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_21;
	cnu_bitSerial_port cnu_converter_port21(
		.serialInOut (cn_serialInOut_21[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_210[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_211[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_212[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_213[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_214[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_215[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_210[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_211[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_212[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_213[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_214[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_215[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_22;
	cnu_bitSerial_port cnu_converter_port22(
		.serialInOut (cn_serialInOut_22[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_220[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_221[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_222[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_223[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_224[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_225[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_220[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_221[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_222[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_223[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_224[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_225[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_23;
	cnu_bitSerial_port cnu_converter_port23(
		.serialInOut (cn_serialInOut_23[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_230[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_231[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_232[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_233[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_234[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_235[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_230[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_231[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_232[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_233[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_234[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_235[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_24;
	cnu_bitSerial_port cnu_converter_port24(
		.serialInOut (cn_serialInOut_24[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_240[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_241[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_242[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_243[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_244[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_245[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_240[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_241[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_242[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_243[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_244[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_245[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_25;
	cnu_bitSerial_port cnu_converter_port25(
		.serialInOut (cn_serialInOut_25[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_250[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_251[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_252[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_253[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_254[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_255[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_250[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_251[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_252[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_253[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_254[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_255[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_26;
	cnu_bitSerial_port cnu_converter_port26(
		.serialInOut (cn_serialInOut_26[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_260[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_261[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_262[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_263[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_264[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_265[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_260[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_261[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_262[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_263[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_264[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_265[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_27;
	cnu_bitSerial_port cnu_converter_port27(
		.serialInOut (cn_serialInOut_27[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_270[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_271[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_272[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_273[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_274[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_275[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_270[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_271[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_272[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_273[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_274[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_275[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_28;
	cnu_bitSerial_port cnu_converter_port28(
		.serialInOut (cn_serialInOut_28[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_280[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_281[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_282[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_283[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_284[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_285[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_280[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_281[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_282[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_283[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_284[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_285[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_29;
	cnu_bitSerial_port cnu_converter_port29(
		.serialInOut (cn_serialInOut_29[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_290[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_291[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_292[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_293[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_294[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_295[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_290[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_291[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_292[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_293[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_294[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_295[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_30;
	cnu_bitSerial_port cnu_converter_port30(
		.serialInOut (cn_serialInOut_30[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_300[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_301[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_302[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_303[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_304[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_305[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_300[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_301[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_302[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_303[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_304[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_305[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_31;
	cnu_bitSerial_port cnu_converter_port31(
		.serialInOut (cn_serialInOut_31[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_310[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_311[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_312[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_313[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_314[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_315[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_310[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_311[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_312[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_313[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_314[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_315[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_32;
	cnu_bitSerial_port cnu_converter_port32(
		.serialInOut (cn_serialInOut_32[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_320[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_321[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_322[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_323[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_324[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_325[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_320[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_321[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_322[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_323[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_324[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_325[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_33;
	cnu_bitSerial_port cnu_converter_port33(
		.serialInOut (cn_serialInOut_33[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_330[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_331[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_332[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_333[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_334[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_335[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_330[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_331[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_332[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_333[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_334[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_335[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_34;
	cnu_bitSerial_port cnu_converter_port34(
		.serialInOut (cn_serialInOut_34[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_340[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_341[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_342[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_343[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_344[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_345[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_340[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_341[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_342[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_343[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_344[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_345[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_35;
	cnu_bitSerial_port cnu_converter_port35(
		.serialInOut (cn_serialInOut_35[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_350[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_351[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_352[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_353[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_354[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_355[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_350[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_351[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_352[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_353[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_354[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_355[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_36;
	cnu_bitSerial_port cnu_converter_port36(
		.serialInOut (cn_serialInOut_36[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_360[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_361[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_362[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_363[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_364[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_365[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_360[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_361[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_362[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_363[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_364[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_365[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_37;
	cnu_bitSerial_port cnu_converter_port37(
		.serialInOut (cn_serialInOut_37[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_370[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_371[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_372[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_373[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_374[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_375[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_370[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_371[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_372[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_373[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_374[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_375[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_38;
	cnu_bitSerial_port cnu_converter_port38(
		.serialInOut (cn_serialInOut_38[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_380[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_381[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_382[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_383[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_384[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_385[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_380[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_381[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_382[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_383[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_384[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_385[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_39;
	cnu_bitSerial_port cnu_converter_port39(
		.serialInOut (cn_serialInOut_39[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_390[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_391[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_392[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_393[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_394[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_395[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_390[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_391[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_392[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_393[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_394[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_395[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_40;
	cnu_bitSerial_port cnu_converter_port40(
		.serialInOut (cn_serialInOut_40[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_400[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_401[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_402[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_403[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_404[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_405[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_400[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_401[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_402[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_403[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_404[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_405[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_41;
	cnu_bitSerial_port cnu_converter_port41(
		.serialInOut (cn_serialInOut_41[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_410[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_411[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_412[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_413[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_414[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_415[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_410[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_411[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_412[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_413[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_414[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_415[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_42;
	cnu_bitSerial_port cnu_converter_port42(
		.serialInOut (cn_serialInOut_42[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_420[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_421[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_422[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_423[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_424[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_425[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_420[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_421[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_422[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_423[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_424[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_425[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_43;
	cnu_bitSerial_port cnu_converter_port43(
		.serialInOut (cn_serialInOut_43[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_430[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_431[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_432[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_433[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_434[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_435[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_430[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_431[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_432[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_433[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_434[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_435[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_44;
	cnu_bitSerial_port cnu_converter_port44(
		.serialInOut (cn_serialInOut_44[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_440[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_441[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_442[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_443[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_444[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_445[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_440[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_441[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_442[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_443[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_444[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_445[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_45;
	cnu_bitSerial_port cnu_converter_port45(
		.serialInOut (cn_serialInOut_45[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_450[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_451[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_452[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_453[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_454[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_455[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_450[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_451[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_452[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_453[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_454[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_455[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_46;
	cnu_bitSerial_port cnu_converter_port46(
		.serialInOut (cn_serialInOut_46[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_460[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_461[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_462[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_463[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_464[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_465[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_460[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_461[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_462[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_463[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_464[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_465[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_47;
	cnu_bitSerial_port cnu_converter_port47(
		.serialInOut (cn_serialInOut_47[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_470[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_471[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_472[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_473[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_474[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_475[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_470[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_471[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_472[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_473[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_474[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_475[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_48;
	cnu_bitSerial_port cnu_converter_port48(
		.serialInOut (cn_serialInOut_48[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_480[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_481[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_482[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_483[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_484[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_485[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_480[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_481[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_482[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_483[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_484[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_485[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_49;
	cnu_bitSerial_port cnu_converter_port49(
		.serialInOut (cn_serialInOut_49[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_490[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_491[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_492[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_493[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_494[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_495[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_490[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_491[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_492[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_493[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_494[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_495[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_50;
	cnu_bitSerial_port cnu_converter_port50(
		.serialInOut (cn_serialInOut_50[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_500[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_501[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_502[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_503[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_504[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_505[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_500[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_501[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_502[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_503[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_504[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_505[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_51;
	cnu_bitSerial_port cnu_converter_port51(
		.serialInOut (cn_serialInOut_51[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_510[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_511[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_512[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_513[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_514[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_515[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_510[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_511[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_512[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_513[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_514[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_515[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_52;
	cnu_bitSerial_port cnu_converter_port52(
		.serialInOut (cn_serialInOut_52[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_520[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_521[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_522[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_523[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_524[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_525[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_520[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_521[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_522[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_523[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_524[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_525[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_53;
	cnu_bitSerial_port cnu_converter_port53(
		.serialInOut (cn_serialInOut_53[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_530[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_531[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_532[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_533[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_534[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_535[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_530[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_531[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_532[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_533[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_534[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_535[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_54;
	cnu_bitSerial_port cnu_converter_port54(
		.serialInOut (cn_serialInOut_54[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_540[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_541[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_542[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_543[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_544[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_545[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_540[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_541[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_542[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_543[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_544[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_545[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_55;
	cnu_bitSerial_port cnu_converter_port55(
		.serialInOut (cn_serialInOut_55[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_550[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_551[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_552[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_553[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_554[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_555[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_550[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_551[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_552[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_553[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_554[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_555[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_56;
	cnu_bitSerial_port cnu_converter_port56(
		.serialInOut (cn_serialInOut_56[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_560[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_561[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_562[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_563[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_564[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_565[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_560[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_561[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_562[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_563[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_564[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_565[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_57;
	cnu_bitSerial_port cnu_converter_port57(
		.serialInOut (cn_serialInOut_57[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_570[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_571[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_572[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_573[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_574[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_575[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_570[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_571[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_572[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_573[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_574[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_575[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_58;
	cnu_bitSerial_port cnu_converter_port58(
		.serialInOut (cn_serialInOut_58[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_580[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_581[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_582[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_583[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_584[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_585[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_580[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_581[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_582[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_583[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_584[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_585[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_59;
	cnu_bitSerial_port cnu_converter_port59(
		.serialInOut (cn_serialInOut_59[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_590[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_591[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_592[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_593[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_594[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_595[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_590[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_591[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_592[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_593[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_594[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_595[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_60;
	cnu_bitSerial_port cnu_converter_port60(
		.serialInOut (cn_serialInOut_60[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_600[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_601[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_602[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_603[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_604[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_605[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_600[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_601[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_602[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_603[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_604[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_605[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_61;
	cnu_bitSerial_port cnu_converter_port61(
		.serialInOut (cn_serialInOut_61[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_610[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_611[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_612[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_613[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_614[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_615[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_610[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_611[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_612[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_613[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_614[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_615[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_62;
	cnu_bitSerial_port cnu_converter_port62(
		.serialInOut (cn_serialInOut_62[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_620[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_621[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_622[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_623[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_624[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_625[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_620[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_621[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_622[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_623[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_624[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_625[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_63;
	cnu_bitSerial_port cnu_converter_port63(
		.serialInOut (cn_serialInOut_63[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_630[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_631[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_632[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_633[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_634[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_635[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_630[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_631[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_632[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_633[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_634[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_635[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_64;
	cnu_bitSerial_port cnu_converter_port64(
		.serialInOut (cn_serialInOut_64[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_640[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_641[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_642[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_643[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_644[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_645[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_640[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_641[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_642[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_643[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_644[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_645[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_65;
	cnu_bitSerial_port cnu_converter_port65(
		.serialInOut (cn_serialInOut_65[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_650[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_651[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_652[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_653[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_654[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_655[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_650[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_651[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_652[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_653[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_654[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_655[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_66;
	cnu_bitSerial_port cnu_converter_port66(
		.serialInOut (cn_serialInOut_66[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_660[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_661[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_662[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_663[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_664[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_665[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_660[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_661[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_662[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_663[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_664[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_665[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_67;
	cnu_bitSerial_port cnu_converter_port67(
		.serialInOut (cn_serialInOut_67[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_670[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_671[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_672[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_673[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_674[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_675[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_670[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_671[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_672[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_673[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_674[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_675[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_68;
	cnu_bitSerial_port cnu_converter_port68(
		.serialInOut (cn_serialInOut_68[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_680[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_681[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_682[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_683[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_684[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_685[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_680[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_681[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_682[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_683[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_684[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_685[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_69;
	cnu_bitSerial_port cnu_converter_port69(
		.serialInOut (cn_serialInOut_69[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_690[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_691[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_692[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_693[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_694[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_695[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_690[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_691[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_692[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_693[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_694[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_695[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_70;
	cnu_bitSerial_port cnu_converter_port70(
		.serialInOut (cn_serialInOut_70[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_700[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_701[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_702[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_703[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_704[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_705[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_700[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_701[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_702[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_703[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_704[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_705[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_71;
	cnu_bitSerial_port cnu_converter_port71(
		.serialInOut (cn_serialInOut_71[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_710[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_711[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_712[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_713[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_714[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_715[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_710[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_711[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_712[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_713[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_714[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_715[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_72;
	cnu_bitSerial_port cnu_converter_port72(
		.serialInOut (cn_serialInOut_72[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_720[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_721[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_722[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_723[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_724[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_725[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_720[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_721[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_722[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_723[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_724[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_725[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_73;
	cnu_bitSerial_port cnu_converter_port73(
		.serialInOut (cn_serialInOut_73[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_730[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_731[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_732[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_733[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_734[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_735[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_730[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_731[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_732[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_733[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_734[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_735[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_74;
	cnu_bitSerial_port cnu_converter_port74(
		.serialInOut (cn_serialInOut_74[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_740[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_741[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_742[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_743[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_744[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_745[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_740[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_741[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_742[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_743[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_744[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_745[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_75;
	cnu_bitSerial_port cnu_converter_port75(
		.serialInOut (cn_serialInOut_75[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_750[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_751[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_752[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_753[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_754[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_755[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_750[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_751[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_752[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_753[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_754[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_755[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_76;
	cnu_bitSerial_port cnu_converter_port76(
		.serialInOut (cn_serialInOut_76[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_760[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_761[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_762[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_763[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_764[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_765[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_760[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_761[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_762[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_763[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_764[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_765[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_77;
	cnu_bitSerial_port cnu_converter_port77(
		.serialInOut (cn_serialInOut_77[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_770[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_771[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_772[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_773[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_774[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_775[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_770[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_771[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_772[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_773[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_774[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_775[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_78;
	cnu_bitSerial_port cnu_converter_port78(
		.serialInOut (cn_serialInOut_78[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_780[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_781[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_782[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_783[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_784[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_785[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_780[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_781[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_782[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_783[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_784[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_785[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_79;
	cnu_bitSerial_port cnu_converter_port79(
		.serialInOut (cn_serialInOut_79[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_790[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_791[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_792[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_793[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_794[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_795[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_790[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_791[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_792[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_793[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_794[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_795[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_80;
	cnu_bitSerial_port cnu_converter_port80(
		.serialInOut (cn_serialInOut_80[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_800[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_801[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_802[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_803[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_804[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_805[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_800[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_801[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_802[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_803[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_804[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_805[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_81;
	cnu_bitSerial_port cnu_converter_port81(
		.serialInOut (cn_serialInOut_81[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_810[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_811[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_812[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_813[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_814[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_815[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_810[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_811[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_812[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_813[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_814[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_815[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_82;
	cnu_bitSerial_port cnu_converter_port82(
		.serialInOut (cn_serialInOut_82[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_820[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_821[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_822[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_823[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_824[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_825[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_820[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_821[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_822[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_823[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_824[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_825[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_83;
	cnu_bitSerial_port cnu_converter_port83(
		.serialInOut (cn_serialInOut_83[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_830[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_831[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_832[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_833[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_834[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_835[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_830[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_831[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_832[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_833[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_834[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_835[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_84;
	cnu_bitSerial_port cnu_converter_port84(
		.serialInOut (cn_serialInOut_84[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_840[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_841[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_842[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_843[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_844[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_845[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_840[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_841[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_842[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_843[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_844[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_845[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_85;
	cnu_bitSerial_port cnu_converter_port85(
		.serialInOut (cn_serialInOut_85[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_850[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_851[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_852[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_853[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_854[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_855[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_850[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_851[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_852[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_853[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_854[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_855[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_86;
	cnu_bitSerial_port cnu_converter_port86(
		.serialInOut (cn_serialInOut_86[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_860[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_861[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_862[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_863[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_864[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_865[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_860[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_861[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_862[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_863[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_864[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_865[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_87;
	cnu_bitSerial_port cnu_converter_port87(
		.serialInOut (cn_serialInOut_87[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_870[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_871[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_872[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_873[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_874[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_875[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_870[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_871[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_872[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_873[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_874[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_875[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_88;
	cnu_bitSerial_port cnu_converter_port88(
		.serialInOut (cn_serialInOut_88[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_880[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_881[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_882[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_883[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_884[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_885[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_880[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_881[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_882[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_883[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_884[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_885[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_89;
	cnu_bitSerial_port cnu_converter_port89(
		.serialInOut (cn_serialInOut_89[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_890[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_891[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_892[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_893[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_894[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_895[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_890[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_891[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_892[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_893[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_894[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_895[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_90;
	cnu_bitSerial_port cnu_converter_port90(
		.serialInOut (cn_serialInOut_90[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_900[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_901[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_902[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_903[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_904[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_905[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_900[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_901[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_902[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_903[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_904[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_905[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_91;
	cnu_bitSerial_port cnu_converter_port91(
		.serialInOut (cn_serialInOut_91[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_910[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_911[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_912[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_913[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_914[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_915[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_910[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_911[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_912[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_913[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_914[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_915[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_92;
	cnu_bitSerial_port cnu_converter_port92(
		.serialInOut (cn_serialInOut_92[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_920[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_921[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_922[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_923[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_924[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_925[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_920[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_921[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_922[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_923[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_924[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_925[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_93;
	cnu_bitSerial_port cnu_converter_port93(
		.serialInOut (cn_serialInOut_93[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_930[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_931[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_932[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_933[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_934[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_935[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_930[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_931[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_932[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_933[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_934[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_935[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_94;
	cnu_bitSerial_port cnu_converter_port94(
		.serialInOut (cn_serialInOut_94[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_940[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_941[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_942[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_943[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_944[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_945[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_940[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_941[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_942[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_943[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_944[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_945[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_95;
	cnu_bitSerial_port cnu_converter_port95(
		.serialInOut (cn_serialInOut_95[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_950[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_951[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_952[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_953[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_954[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_955[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_950[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_951[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_952[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_953[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_954[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_955[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_96;
	cnu_bitSerial_port cnu_converter_port96(
		.serialInOut (cn_serialInOut_96[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_960[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_961[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_962[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_963[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_964[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_965[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_960[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_961[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_962[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_963[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_964[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_965[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_97;
	cnu_bitSerial_port cnu_converter_port97(
		.serialInOut (cn_serialInOut_97[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_970[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_971[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_972[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_973[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_974[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_975[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_970[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_971[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_972[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_973[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_974[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_975[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_98;
	cnu_bitSerial_port cnu_converter_port98(
		.serialInOut (cn_serialInOut_98[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_980[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_981[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_982[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_983[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_984[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_985[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_980[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_981[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_982[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_983[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_984[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_985[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_99;
	cnu_bitSerial_port cnu_converter_port99(
		.serialInOut (cn_serialInOut_99[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_990[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_991[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_992[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_993[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_994[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_995[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_990[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_991[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_992[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_993[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_994[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_995[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_100;
	cnu_bitSerial_port cnu_converter_port100(
		.serialInOut (cn_serialInOut_100[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_1000[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_1001[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_1002[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_1003[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_1004[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_1005[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_1000[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_1001[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_1002[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_1003[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_1004[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_1005[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	wire [`CN_DEGREE-1:0] cn_serialInOut_101;
	cnu_bitSerial_port cnu_converter_port101(
		.serialInOut (cn_serialInOut_101[`CN_DEGREE-1:0]),
		.v2c_parallelOut_0 (v2c_parallelOut_1010[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_1 (v2c_parallelOut_1011[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_2 (v2c_parallelOut_1012[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_3 (v2c_parallelOut_1013[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_4 (v2c_parallelOut_1014[`DATAPATH_WIDTH-1:0]),
		.v2c_parallelOut_5 (v2c_parallelOut_1015[`DATAPATH_WIDTH-1:0]),
		
		.c2v_parallelIn_0 (c2v_parallelIn_1010[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_1 (c2v_parallelIn_1011[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_2 (c2v_parallelIn_1012[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_3 (c2v_parallelIn_1013[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_4 (c2v_parallelIn_1014[`DATAPATH_WIDTH-1:0]),
		.c2v_parallelIn_5 (c2v_parallelIn_1015[`DATAPATH_WIDTH-1:0]),
		.load (load[0]),
		.parallel_en (parallel_en[0]),
		.serial_clk (serial_clk)
	);
	
	vnu_bitSerial_port vnu_converter_port0 (
		.serialInOut ({cn_serialInOut_72[0], cn_serialInOut_83[0], cn_serialInOut_80[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port1 (
		.serialInOut ({cn_serialInOut_62[0], cn_serialInOut_44[0], cn_serialInOut_25[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port2 (
		.serialInOut ({cn_serialInOut_16[0], cn_serialInOut_76[0], cn_serialInOut_54[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port3 (
		.serialInOut ({cn_serialInOut_73[0], cn_serialInOut_46[0], cn_serialInOut_23[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port4 (
		.serialInOut ({cn_serialInOut_8[0], cn_serialInOut_9[0], cn_serialInOut_51[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port5 (
		.serialInOut ({cn_serialInOut_61[0], cn_serialInOut_62[1], cn_serialInOut_43[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port6 (
		.serialInOut ({cn_serialInOut_37[0], cn_serialInOut_38[0], cn_serialInOut_34[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port7 (
		.serialInOut ({cn_serialInOut_59[0], cn_serialInOut_3[0], cn_serialInOut_99[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port8 (
		.serialInOut ({cn_serialInOut_81[0], cn_serialInOut_97[0], cn_serialInOut_62[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port9 (
		.serialInOut ({cn_serialInOut_39[0], cn_serialInOut_79[0], cn_serialInOut_67[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port10 (
		.serialInOut ({cn_serialInOut_90[0], cn_serialInOut_80[1], cn_serialInOut_17[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port11 (
		.serialInOut ({cn_serialInOut_85[0], cn_serialInOut_87[0], cn_serialInOut_98[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port12 (
		.serialInOut ({cn_serialInOut_76[1], cn_serialInOut_70[0], cn_serialInOut_64[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port13 (
		.serialInOut ({cn_serialInOut_28[0], cn_serialInOut_8[1], cn_serialInOut_32[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port14 (
		.serialInOut ({cn_serialInOut_14[0], cn_serialInOut_40[0], cn_serialInOut_33[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port15 (
		.serialInOut ({cn_serialInOut_74[0], cn_serialInOut_10[0], cn_serialInOut_21[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port16 (
		.serialInOut ({cn_serialInOut_47[0], cn_serialInOut_23[1], cn_serialInOut_94[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port17 (
		.serialInOut ({cn_serialInOut_21[1], cn_serialInOut_43[1], cn_serialInOut_59[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port18 (
		.serialInOut ({cn_serialInOut_4[0], cn_serialInOut_18[0], cn_serialInOut_40[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port19 (
		.serialInOut ({cn_serialInOut_30[0], cn_serialInOut_21[2], cn_serialInOut_42[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port20 (
		.serialInOut ({cn_serialInOut_20[0], cn_serialInOut_17[1], cn_serialInOut_55[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port21 (
		.serialInOut ({cn_serialInOut_82[0], cn_serialInOut_50[0], cn_serialInOut_48[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port22 (
		.serialInOut ({cn_serialInOut_78[0], cn_serialInOut_6[0], cn_serialInOut_87[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port23 (
		.serialInOut ({cn_serialInOut_35[0], cn_serialInOut_66[0], cn_serialInOut_4[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port24 (
		.serialInOut ({cn_serialInOut_83[1], cn_serialInOut_74[1], cn_serialInOut_31[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port25 (
		.serialInOut ({cn_serialInOut_0[0], cn_serialInOut_78[1], cn_serialInOut_37[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port26 (
		.serialInOut ({cn_serialInOut_42[1], cn_serialInOut_81[1], cn_serialInOut_74[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port27 (
		.serialInOut ({cn_serialInOut_1[0], cn_serialInOut_0[1], cn_serialInOut_22[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port28 (
		.serialInOut ({cn_serialInOut_32[1], cn_serialInOut_60[0], cn_serialInOut_82[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port29 (
		.serialInOut ({cn_serialInOut_68[0], cn_serialInOut_2[0], cn_serialInOut_29[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port30 (
		.serialInOut ({cn_serialInOut_27[0], cn_serialInOut_4[2], cn_serialInOut_76[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port31 (
		.serialInOut ({cn_serialInOut_7[0], cn_serialInOut_55[1], cn_serialInOut_3[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port32 (
		.serialInOut ({cn_serialInOut_52[0], cn_serialInOut_75[0], cn_serialInOut_35[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port33 (
		.serialInOut ({cn_serialInOut_95[0], cn_serialInOut_27[1], cn_serialInOut_101[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port34 (
		.serialInOut ({cn_serialInOut_43[2], cn_serialInOut_16[1], cn_serialInOut_47[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port35 (
		.serialInOut ({cn_serialInOut_91[0], cn_serialInOut_25[1], cn_serialInOut_73[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port36 (
		.serialInOut ({cn_serialInOut_55[2], cn_serialInOut_68[1], cn_serialInOut_10[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port37 (
		.serialInOut ({cn_serialInOut_17[2], cn_serialInOut_67[1], cn_serialInOut_49[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port38 (
		.serialInOut ({cn_serialInOut_71[0], cn_serialInOut_33[1], cn_serialInOut_36[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port39 (
		.serialInOut ({cn_serialInOut_24[0], cn_serialInOut_36[1], cn_serialInOut_75[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port40 (
		.serialInOut ({cn_serialInOut_22[1], cn_serialInOut_29[1], cn_serialInOut_20[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port41 (
		.serialInOut ({cn_serialInOut_6[1], cn_serialInOut_28[1], cn_serialInOut_39[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port42 (
		.serialInOut ({cn_serialInOut_70[1], cn_serialInOut_77[0], cn_serialInOut_38[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port43 (
		.serialInOut ({cn_serialInOut_12[0], cn_serialInOut_1[1], cn_serialInOut_95[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port44 (
		.serialInOut ({cn_serialInOut_54[1], cn_serialInOut_32[2], cn_serialInOut_50[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port45 (
		.serialInOut ({cn_serialInOut_48[1], cn_serialInOut_63[0], cn_serialInOut_15[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port46 (
		.serialInOut ({cn_serialInOut_36[2], cn_serialInOut_65[0], cn_serialInOut_53[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port47 (
		.serialInOut ({cn_serialInOut_49[1], cn_serialInOut_35[2], cn_serialInOut_88[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port48 (
		.serialInOut ({cn_serialInOut_44[1], cn_serialInOut_14[1], cn_serialInOut_56[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port49 (
		.serialInOut ({cn_serialInOut_87[2], cn_serialInOut_34[1], cn_serialInOut_14[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port50 (
		.serialInOut ({cn_serialInOut_56[1], cn_serialInOut_101[1], cn_serialInOut_77[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port51 (
		.serialInOut ({cn_serialInOut_97[1], cn_serialInOut_26[0], cn_serialInOut_70[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port52 (
		.serialInOut ({cn_serialInOut_26[1], cn_serialInOut_51[1], cn_serialInOut_93[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port53 (
		.serialInOut ({cn_serialInOut_67[2], cn_serialInOut_19[0], cn_serialInOut_86[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port54 (
		.serialInOut ({cn_serialInOut_88[1], cn_serialInOut_37[2], cn_serialInOut_7[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port55 (
		.serialInOut ({cn_serialInOut_23[2], cn_serialInOut_93[1], cn_serialInOut_52[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port56 (
		.serialInOut ({cn_serialInOut_10[2], cn_serialInOut_49[2], cn_serialInOut_18[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port57 (
		.serialInOut ({cn_serialInOut_13[0], cn_serialInOut_82[2], cn_serialInOut_97[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port58 (
		.serialInOut ({cn_serialInOut_75[2], cn_serialInOut_54[2], cn_serialInOut_1[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port59 (
		.serialInOut ({cn_serialInOut_40[2], cn_serialInOut_69[0], cn_serialInOut_61[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port60 (
		.serialInOut ({cn_serialInOut_77[2], cn_serialInOut_85[1], cn_serialInOut_13[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port61 (
		.serialInOut ({cn_serialInOut_2[1], cn_serialInOut_20[2], cn_serialInOut_58[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port62 (
		.serialInOut ({cn_serialInOut_63[1], cn_serialInOut_22[2], cn_serialInOut_45[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port63 (
		.serialInOut ({cn_serialInOut_46[1], cn_serialInOut_42[2], cn_serialInOut_44[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port64 (
		.serialInOut ({cn_serialInOut_94[1], cn_serialInOut_30[1], cn_serialInOut_0[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port65 (
		.serialInOut ({cn_serialInOut_84[0], cn_serialInOut_58[1], cn_serialInOut_83[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port66 (
		.serialInOut ({cn_serialInOut_93[2], cn_serialInOut_53[1], cn_serialInOut_100[0]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port67 (
		.serialInOut ({cn_serialInOut_92[0], cn_serialInOut_5[0], cn_serialInOut_30[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port68 (
		.serialInOut ({cn_serialInOut_58[2], cn_serialInOut_94[2], cn_serialInOut_60[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port69 (
		.serialInOut ({cn_serialInOut_57[0], cn_serialInOut_72[1], cn_serialInOut_46[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port70 (
		.serialInOut ({cn_serialInOut_53[2], cn_serialInOut_86[1], cn_serialInOut_6[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port71 (
		.serialInOut ({cn_serialInOut_51[2], cn_serialInOut_96[0], cn_serialInOut_78[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port72 (
		.serialInOut ({cn_serialInOut_11[0], cn_serialInOut_89[0], cn_serialInOut_27[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port73 (
		.serialInOut ({cn_serialInOut_29[2], cn_serialInOut_98[1], cn_serialInOut_96[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port74 (
		.serialInOut ({cn_serialInOut_41[0], cn_serialInOut_99[1], cn_serialInOut_72[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port75 (
		.serialInOut ({cn_serialInOut_100[1], cn_serialInOut_61[2], cn_serialInOut_19[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port76 (
		.serialInOut ({cn_serialInOut_79[1], cn_serialInOut_95[2], cn_serialInOut_84[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port77 (
		.serialInOut ({cn_serialInOut_99[2], cn_serialInOut_57[1], cn_serialInOut_90[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port78 (
		.serialInOut ({cn_serialInOut_18[2], cn_serialInOut_15[1], cn_serialInOut_5[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port79 (
		.serialInOut ({cn_serialInOut_98[2], cn_serialInOut_48[2], cn_serialInOut_71[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port80 (
		.serialInOut ({cn_serialInOut_69[1], cn_serialInOut_91[1], cn_serialInOut_16[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port81 (
		.serialInOut ({cn_serialInOut_89[1], cn_serialInOut_92[1], cn_serialInOut_68[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port82 (
		.serialInOut ({cn_serialInOut_9[1], cn_serialInOut_39[2], cn_serialInOut_24[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port83 (
		.serialInOut ({cn_serialInOut_38[2], cn_serialInOut_71[2], cn_serialInOut_81[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port84 (
		.serialInOut ({cn_serialInOut_66[1], cn_serialInOut_73[2], cn_serialInOut_11[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port85 (
		.serialInOut ({cn_serialInOut_3[2], cn_serialInOut_64[1], cn_serialInOut_26[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port86 (
		.serialInOut ({cn_serialInOut_19[2], cn_serialInOut_84[2], cn_serialInOut_89[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port87 (
		.serialInOut ({cn_serialInOut_101[2], cn_serialInOut_12[1], cn_serialInOut_91[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port88 (
		.serialInOut ({cn_serialInOut_45[1], cn_serialInOut_7[2], cn_serialInOut_8[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port89 (
		.serialInOut ({cn_serialInOut_34[2], cn_serialInOut_45[2], cn_serialInOut_9[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port90 (
		.serialInOut ({cn_serialInOut_96[2], cn_serialInOut_52[2], cn_serialInOut_92[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port91 (
		.serialInOut ({cn_serialInOut_65[1], cn_serialInOut_47[2], cn_serialInOut_41[1]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port92 (
		.serialInOut ({cn_serialInOut_86[2], cn_serialInOut_88[2], cn_serialInOut_63[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port93 (
		.serialInOut ({cn_serialInOut_25[2], cn_serialInOut_24[2], cn_serialInOut_57[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port94 (
		.serialInOut ({cn_serialInOut_5[2], cn_serialInOut_56[2], cn_serialInOut_66[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port95 (
		.serialInOut ({cn_serialInOut_64[2], cn_serialInOut_11[2], cn_serialInOut_2[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port96 (
		.serialInOut ({cn_serialInOut_60[2], cn_serialInOut_90[2], cn_serialInOut_65[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port97 (
		.serialInOut ({cn_serialInOut_80[2], cn_serialInOut_100[2], cn_serialInOut_28[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port98 (
		.serialInOut ({cn_serialInOut_50[2], cn_serialInOut_59[2], cn_serialInOut_85[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port99 (
		.serialInOut ({cn_serialInOut_15[2], cn_serialInOut_13[2], cn_serialInOut_79[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port100 (
		.serialInOut ({cn_serialInOut_33[2], cn_serialInOut_31[1], cn_serialInOut_69[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port101 (
		.serialInOut ({cn_serialInOut_31[2], cn_serialInOut_41[2], cn_serialInOut_12[2]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port102 (
		.serialInOut ({cn_serialInOut_71[3], cn_serialInOut_16[3], cn_serialInOut_44[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port103 (
		.serialInOut ({cn_serialInOut_51[3], cn_serialInOut_13[3], cn_serialInOut_21[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port104 (
		.serialInOut ({cn_serialInOut_48[3], cn_serialInOut_52[3], cn_serialInOut_1[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port105 (
		.serialInOut ({cn_serialInOut_94[3], cn_serialInOut_75[3], cn_serialInOut_59[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port106 (
		.serialInOut ({cn_serialInOut_38[3], cn_serialInOut_56[3], cn_serialInOut_25[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port107 (
		.serialInOut ({cn_serialInOut_31[3], cn_serialInOut_59[4], cn_serialInOut_47[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port108 (
		.serialInOut ({cn_serialInOut_1[4], cn_serialInOut_77[3], cn_serialInOut_7[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port109 (
		.serialInOut ({cn_serialInOut_91[3], cn_serialInOut_2[3], cn_serialInOut_53[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port110 (
		.serialInOut ({cn_serialInOut_70[3], cn_serialInOut_54[3], cn_serialInOut_41[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port111 (
		.serialInOut ({cn_serialInOut_22[3], cn_serialInOut_4[3], cn_serialInOut_61[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port112 (
		.serialInOut ({cn_serialInOut_34[3], cn_serialInOut_98[3], cn_serialInOut_49[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port113 (
		.serialInOut ({cn_serialInOut_36[3], cn_serialInOut_30[3], cn_serialInOut_17[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port114 (
		.serialInOut ({cn_serialInOut_23[3], cn_serialInOut_83[3], cn_serialInOut_11[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port115 (
		.serialInOut ({cn_serialInOut_13[4], cn_serialInOut_96[3], cn_serialInOut_55[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port116 (
		.serialInOut ({cn_serialInOut_93[3], cn_serialInOut_39[3], cn_serialInOut_43[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port117 (
		.serialInOut ({cn_serialInOut_21[4], cn_serialInOut_73[3], cn_serialInOut_62[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port118 (
		.serialInOut ({cn_serialInOut_62[4], cn_serialInOut_48[4], cn_serialInOut_27[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port119 (
		.serialInOut ({cn_serialInOut_41[4], cn_serialInOut_95[3], cn_serialInOut_77[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port120 (
		.serialInOut ({cn_serialInOut_100[3], cn_serialInOut_26[3], cn_serialInOut_84[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port121 (
		.serialInOut ({cn_serialInOut_54[4], cn_serialInOut_74[3], cn_serialInOut_98[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port122 (
		.serialInOut ({cn_serialInOut_39[4], cn_serialInOut_8[3], cn_serialInOut_66[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port123 (
		.serialInOut ({cn_serialInOut_60[3], cn_serialInOut_27[4], cn_serialInOut_96[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port124 (
		.serialInOut ({cn_serialInOut_75[4], cn_serialInOut_100[4], cn_serialInOut_15[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port125 (
		.serialInOut ({cn_serialInOut_87[3], cn_serialInOut_94[4], cn_serialInOut_32[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port126 (
		.serialInOut ({cn_serialInOut_4[4], cn_serialInOut_32[4], cn_serialInOut_36[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port127 (
		.serialInOut ({cn_serialInOut_67[3], cn_serialInOut_60[4], cn_serialInOut_26[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port128 (
		.serialInOut ({cn_serialInOut_64[3], cn_serialInOut_51[4], cn_serialInOut_37[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port129 (
		.serialInOut ({cn_serialInOut_19[3], cn_serialInOut_41[5], cn_serialInOut_14[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port130 (
		.serialInOut ({cn_serialInOut_59[5], cn_serialInOut_22[4], cn_serialInOut_83[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port131 (
		.serialInOut ({cn_serialInOut_66[4], cn_serialInOut_72[3], cn_serialInOut_51[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port132 (
		.serialInOut ({cn_serialInOut_24[3], cn_serialInOut_65[3], cn_serialInOut_52[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port133 (
		.serialInOut ({cn_serialInOut_50[3], cn_serialInOut_76[3], cn_serialInOut_20[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port134 (
		.serialInOut ({cn_serialInOut_80[3], cn_serialInOut_61[4], cn_serialInOut_0[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port135 (
		.serialInOut ({cn_serialInOut_65[4], cn_serialInOut_20[4], cn_serialInOut_95[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port136 (
		.serialInOut ({cn_serialInOut_74[4], cn_serialInOut_55[4], cn_serialInOut_82[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port137 (
		.serialInOut ({cn_serialInOut_7[4], cn_serialInOut_12[3], cn_serialInOut_18[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port138 (
		.serialInOut ({cn_serialInOut_29[3], cn_serialInOut_18[4], cn_serialInOut_50[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port139 (
		.serialInOut ({cn_serialInOut_101[3], cn_serialInOut_89[3], cn_serialInOut_57[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port140 (
		.serialInOut ({cn_serialInOut_96[5], cn_serialInOut_10[3], cn_serialInOut_67[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port141 (
		.serialInOut ({cn_serialInOut_88[3], cn_serialInOut_14[4], cn_serialInOut_97[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port142 (
		.serialInOut ({cn_serialInOut_43[4], cn_serialInOut_19[4], cn_serialInOut_34[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port143 (
		.serialInOut ({cn_serialInOut_73[4], cn_serialInOut_34[5], cn_serialInOut_4[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port144 (
		.serialInOut ({cn_serialInOut_25[4], cn_serialInOut_71[4], cn_serialInOut_58[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port145 (
		.serialInOut ({cn_serialInOut_9[3], cn_serialInOut_87[4], cn_serialInOut_93[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port146 (
		.serialInOut ({cn_serialInOut_45[3], cn_serialInOut_68[3], cn_serialInOut_99[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port147 (
		.serialInOut ({cn_serialInOut_15[4], cn_serialInOut_53[4], cn_serialInOut_76[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port148 (
		.serialInOut ({cn_serialInOut_90[3], cn_serialInOut_5[3], cn_serialInOut_73[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port149 (
		.serialInOut ({cn_serialInOut_12[4], cn_serialInOut_63[3], cn_serialInOut_100[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port150 (
		.serialInOut ({cn_serialInOut_46[3], cn_serialInOut_31[4], cn_serialInOut_39[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port151 (
		.serialInOut ({cn_serialInOut_49[4], cn_serialInOut_23[4], cn_serialInOut_89[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port152 (
		.serialInOut ({cn_serialInOut_37[4], cn_serialInOut_47[4], cn_serialInOut_45[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port153 (
		.serialInOut ({cn_serialInOut_85[3], cn_serialInOut_84[4], cn_serialInOut_46[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port154 (
		.serialInOut ({cn_serialInOut_5[4], cn_serialInOut_50[5], cn_serialInOut_33[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port155 (
		.serialInOut ({cn_serialInOut_6[3], cn_serialInOut_67[5], cn_serialInOut_35[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port156 (
		.serialInOut ({cn_serialInOut_55[5], cn_serialInOut_6[4], cn_serialInOut_30[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port157 (
		.serialInOut ({cn_serialInOut_68[4], cn_serialInOut_91[4], cn_serialInOut_60[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port158 (
		.serialInOut ({cn_serialInOut_47[5], cn_serialInOut_38[4], cn_serialInOut_42[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port159 (
		.serialInOut ({cn_serialInOut_30[5], cn_serialInOut_70[4], cn_serialInOut_63[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port160 (
		.serialInOut ({cn_serialInOut_32[5], cn_serialInOut_7[5], cn_serialInOut_92[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port161 (
		.serialInOut ({cn_serialInOut_78[3], cn_serialInOut_3[3], cn_serialInOut_16[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port162 (
		.serialInOut ({cn_serialInOut_97[4], cn_serialInOut_36[5], cn_serialInOut_94[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port163 (
		.serialInOut ({cn_serialInOut_76[5], cn_serialInOut_86[3], cn_serialInOut_24[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port164 (
		.serialInOut ({cn_serialInOut_18[5], cn_serialInOut_66[5], cn_serialInOut_48[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port165 (
		.serialInOut ({cn_serialInOut_86[4], cn_serialInOut_1[5], cn_serialInOut_68[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port166 (
		.serialInOut ({cn_serialInOut_0[4], cn_serialInOut_21[5], cn_serialInOut_9[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port167 (
		.serialInOut ({cn_serialInOut_63[5], cn_serialInOut_28[3], cn_serialInOut_87[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port168 (
		.serialInOut ({cn_serialInOut_69[3], cn_serialInOut_90[4], cn_serialInOut_64[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port169 (
		.serialInOut ({cn_serialInOut_83[5], cn_serialInOut_24[5], cn_serialInOut_101[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port170 (
		.serialInOut ({cn_serialInOut_98[5], cn_serialInOut_44[4], cn_serialInOut_65[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port171 (
		.serialInOut ({cn_serialInOut_57[4], cn_serialInOut_17[4], cn_serialInOut_56[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port172 (
		.serialInOut ({cn_serialInOut_3[4], cn_serialInOut_0[5], cn_serialInOut_69[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port173 (
		.serialInOut ({cn_serialInOut_11[4], cn_serialInOut_29[4], cn_serialInOut_71[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port174 (
		.serialInOut ({cn_serialInOut_81[3], cn_serialInOut_88[4], cn_serialInOut_31[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port175 (
		.serialInOut ({cn_serialInOut_14[5], cn_serialInOut_46[5], cn_serialInOut_54[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port176 (
		.serialInOut ({cn_serialInOut_17[5], cn_serialInOut_58[4], cn_serialInOut_23[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port177 (
		.serialInOut ({cn_serialInOut_20[5], cn_serialInOut_80[4], cn_serialInOut_12[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port178 (
		.serialInOut ({cn_serialInOut_53[5], cn_serialInOut_99[4], cn_serialInOut_28[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port179 (
		.serialInOut ({cn_serialInOut_56[5], cn_serialInOut_49[5], cn_serialInOut_3[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port180 (
		.serialInOut ({cn_serialInOut_89[5], cn_serialInOut_93[5], cn_serialInOut_22[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port181 (
		.serialInOut ({cn_serialInOut_33[4], cn_serialInOut_9[5], cn_serialInOut_78[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port182 (
		.serialInOut ({cn_serialInOut_92[4], cn_serialInOut_43[5], cn_serialInOut_88[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port183 (
		.serialInOut ({cn_serialInOut_72[4], cn_serialInOut_101[5], cn_serialInOut_40[3]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port184 (
		.serialInOut ({cn_serialInOut_79[3], cn_serialInOut_25[5], cn_serialInOut_81[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port185 (
		.serialInOut ({cn_serialInOut_10[4], cn_serialInOut_64[5], cn_serialInOut_91[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port186 (
		.serialInOut ({cn_serialInOut_44[5], cn_serialInOut_40[4], cn_serialInOut_86[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port187 (
		.serialInOut ({cn_serialInOut_27[5], cn_serialInOut_82[4], cn_serialInOut_70[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port188 (
		.serialInOut ({cn_serialInOut_84[5], cn_serialInOut_33[5], cn_serialInOut_38[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port189 (
		.serialInOut ({cn_serialInOut_8[4], cn_serialInOut_81[5], cn_serialInOut_13[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port190 (
		.serialInOut ({cn_serialInOut_2[4], cn_serialInOut_35[4], cn_serialInOut_19[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port191 (
		.serialInOut ({cn_serialInOut_82[5], cn_serialInOut_85[4], cn_serialInOut_75[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port192 (
		.serialInOut ({cn_serialInOut_28[5], cn_serialInOut_69[5], cn_serialInOut_79[4]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port193 (
		.serialInOut ({cn_serialInOut_42[4], cn_serialInOut_11[5], cn_serialInOut_8[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port194 (
		.serialInOut ({cn_serialInOut_77[5], cn_serialInOut_62[5], cn_serialInOut_72[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port195 (
		.serialInOut ({cn_serialInOut_26[5], cn_serialInOut_45[5], cn_serialInOut_29[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port196 (
		.serialInOut ({cn_serialInOut_58[5], cn_serialInOut_15[5], cn_serialInOut_85[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port197 (
		.serialInOut ({cn_serialInOut_61[5], cn_serialInOut_57[5], cn_serialInOut_5[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port198 (
		.serialInOut ({cn_serialInOut_40[5], cn_serialInOut_97[5], cn_serialInOut_90[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port199 (
		.serialInOut ({cn_serialInOut_95[5], cn_serialInOut_92[5], cn_serialInOut_10[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port200 (
		.serialInOut ({cn_serialInOut_52[5], cn_serialInOut_42[5], cn_serialInOut_80[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port201 (
		.serialInOut ({cn_serialInOut_35[5], cn_serialInOut_78[5], cn_serialInOut_74[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port202 (
		.serialInOut ({cn_serialInOut_16[5], cn_serialInOut_37[5], cn_serialInOut_2[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);

	vnu_bitSerial_port vnu_converter_port203 (
		.serialInOut ({cn_serialInOut_99[5], cn_serialInOut_79[5], cn_serialInOut_6[5]}),
		.load (load[1]),
		.parallel_en (parallel_en[1]),
		.serial_clk (serial_clk)
	);
endmodule