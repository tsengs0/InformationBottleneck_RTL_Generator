`include "define.v"

module ib_lut_cnu_f0 (
	output reg [`QUAN_SIZE-1:0] t_c,
	
	input wire [`QUAN_SIZE-1:0] y0,
	input wire [`QUAN_SIZE-1:0] y1
);
always @(y0, y1) begin
	case({y0, y1}) 
		{`QUAN_SIZE'd0, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd15;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd14;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd1;
		{`QUAN_SIZE'd0, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd0;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd14;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd14;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd1;
		{`QUAN_SIZE'd1, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd1;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd2, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd3, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd4, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd5, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd6, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd7, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd8, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd9, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd10, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd11, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd12, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd13, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd1;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd1;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd14;
		{`QUAN_SIZE'd14, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd14;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd0}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd0;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd1}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd1;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd2}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd2;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd3}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd3;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd4}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd4;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd5}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd5;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd6}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd6;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd7}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd7;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd8}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd8;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd9}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd9;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd10}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd10;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd11}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd11;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd12}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd12;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd13}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd13;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd14}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd14;
		{`QUAN_SIZE'd15, `QUAN_SIZE'd15}: t_c[`QUAN_SIZE-1:0] <= `QUAN_SIZE'd15;
	endcase
end

endmodule 
