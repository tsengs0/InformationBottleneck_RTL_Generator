`include "define.vh"

`ifdef SCHED_4_6
module mem_subsystem_top_submatrix_9 #(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 85,
	parameter LAYER_NUM = 3,
	parameter CH_DATA_WIDTH = CHECK_PARALLELISM*QUAN_SIZE,
	// Parameters of extrinsic RAMs
	parameter RAM_PORTA_RANGE = 9, // 9 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port A,
	parameter RAM_PORTB_RANGE = 9, // 8 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port b, 
	parameter MEM_DEVICE_NUM = 9,
	parameter DEPTH = 1024,
	parameter DATA_WIDTH = 36,
	parameter FRAG_DATA_WIDTH = 16,
	parameter ADDR_WIDTH = $clog2(DEPTH)
) (
	output wire [CHECK_PARALLELISM-1:0] vnu_pa_msg_bit0,
	output wire [CH_DATA_WIDTH-1:0] pa_to_ch_ram,
	// The memory Dout port to variable nodes as instrinsic messages
	output wire [QUAN_SIZE-1:0] mem_to_vnu_0,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_1,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_2,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_3,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_4,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_5,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_6,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_7,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_8,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_9,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_10,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_11,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_12,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_13,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_14,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_15,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_16,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_17,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_18,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_19,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_20,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_21,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_22,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_23,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_24,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_25,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_26,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_27,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_28,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_29,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_30,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_31,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_32,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_33,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_34,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_35,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_36,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_37,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_38,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_39,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_40,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_41,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_42,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_43,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_44,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_45,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_46,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_47,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_48,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_49,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_50,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_51,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_52,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_53,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_54,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_55,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_56,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_57,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_58,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_59,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_60,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_61,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_62,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_63,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_64,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_65,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_66,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_67,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_68,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_69,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_70,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_71,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_72,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_73,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_74,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_75,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_76,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_77,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_78,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_79,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_80,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_81,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_82,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_83,
	output wire [QUAN_SIZE-1:0] mem_to_vnu_84,
	// The memory Dout port to check nodes as instrinsic messages
	output wire [QUAN_SIZE-1:0] mem_to_cnu_0,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_1,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_2,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_3,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_4,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_5,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_6,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_7,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_8,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_9,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_10,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_11,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_12,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_13,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_14,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_15,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_16,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_17,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_18,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_19,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_20,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_21,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_22,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_23,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_24,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_25,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_26,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_27,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_28,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_29,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_30,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_31,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_32,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_33,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_34,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_35,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_36,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_37,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_38,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_39,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_40,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_41,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_42,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_43,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_44,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_45,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_46,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_47,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_48,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_49,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_50,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_51,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_52,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_53,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_54,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_55,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_56,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_57,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_58,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_59,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_60,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_61,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_62,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_63,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_64,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_65,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_66,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_67,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_68,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_69,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_70,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_71,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_72,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_73,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_74,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_75,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_76,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_77,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_78,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_79,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_80,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_81,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_82,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_83,
	output wire [QUAN_SIZE-1:0] mem_to_cnu_84,
	// The varible extrinsic message written back onto memory through BS and PA
	input wire [QUAN_SIZE-1:0] vnu_to_mem_0,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_1,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_2,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_3,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_4,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_5,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_6,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_7,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_8,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_9,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_10,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_11,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_12,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_13,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_14,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_15,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_16,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_17,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_18,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_19,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_20,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_21,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_22,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_23,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_24,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_25,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_26,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_27,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_28,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_29,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_30,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_31,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_32,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_33,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_34,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_35,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_36,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_37,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_38,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_39,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_40,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_41,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_42,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_43,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_44,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_45,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_46,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_47,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_48,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_49,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_50,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_51,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_52,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_53,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_54,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_55,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_56,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_57,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_58,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_59,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_60,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_61,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_62,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_63,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_64,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_65,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_66,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_67,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_68,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_69,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_70,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_71,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_72,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_73,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_74,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_75,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_76,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_77,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_78,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_79,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_80,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_81,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_82,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_83,
	input wire [QUAN_SIZE-1:0] vnu_to_mem_84,
	// The check extrinsic message written back onto memory through BS and PA
	input wire [QUAN_SIZE-1:0] cnu_to_mem_0,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_1,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_2,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_3,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_4,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_5,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_6,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_7,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_8,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_9,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_10,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_11,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_12,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_13,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_14,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_15,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_16,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_17,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_18,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_19,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_20,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_21,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_22,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_23,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_24,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_25,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_26,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_27,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_28,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_29,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_30,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_31,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_32,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_33,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_34,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_35,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_36,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_37,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_38,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_39,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_40,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_41,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_42,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_43,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_44,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_45,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_46,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_47,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_48,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_49,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_50,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_51,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_52,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_53,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_54,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_55,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_56,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_57,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_58,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_59,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_60,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_61,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_62,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_63,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_64,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_65,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_66,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_67,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_68,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_69,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_70,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_71,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_72,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_73,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_74,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_75,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_76,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_77,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_78,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_79,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_80,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_81,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_82,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_83,
	input wire [QUAN_SIZE-1:0] cnu_to_mem_84,

	input wire [ADDR_WIDTH-1:0] cnu_sync_addr,
	input wire [ADDR_WIDTH-1:0] vnu_sync_addr,
	input wire [LAYER_NUM-1:0] cnu_layer_status,
	input wire [LAYER_NUM-1:0] vnu_layer_status,
	input wire [1:0] last_row_chunk, // [0]: check; [1]: variable
	input wire [1:0] we, // [0]: check; [1]: variable
	input wire sys_clk,
	input wire rstn
);

/*-------------------------------------------------------*/
// Page alignment of Check nodes
wire [QUAN_SIZE-1:0] cnu_pa_msg [CHECK_PARALLELISM-1:0];
ram_pageAlign_interface_submatrix_9 #(
	.QUAN_SIZE(QUAN_SIZE),
	.CHECK_PARALLELISM(CHECK_PARALLELISM),
	.LAYER_NUM(LAYER_NUM)
) cnu_ram_pageAlign_interface_submatrix_9 (
	.msg_out_0       (cnu_pa_msg[0 ]),
	.msg_out_1       (cnu_pa_msg[1 ]),
	.msg_out_2       (cnu_pa_msg[2 ]),
	.msg_out_3       (cnu_pa_msg[3 ]),
	.msg_out_4       (cnu_pa_msg[4 ]),
	.msg_out_5       (cnu_pa_msg[5 ]),
	.msg_out_6       (cnu_pa_msg[6 ]),
	.msg_out_7       (cnu_pa_msg[7 ]),
	.msg_out_8       (cnu_pa_msg[8 ]),
	.msg_out_9       (cnu_pa_msg[9 ]),
	.msg_out_10      (cnu_pa_msg[10]),
	.msg_out_11      (cnu_pa_msg[11]),
	.msg_out_12      (cnu_pa_msg[12]),
	.msg_out_13      (cnu_pa_msg[13]),
	.msg_out_14      (cnu_pa_msg[14]),
	.msg_out_15      (cnu_pa_msg[15]),
	.msg_out_16      (cnu_pa_msg[16]),
	.msg_out_17      (cnu_pa_msg[17]),
	.msg_out_18      (cnu_pa_msg[18]),
	.msg_out_19      (cnu_pa_msg[19]),
	.msg_out_20      (cnu_pa_msg[20]),
	.msg_out_21      (cnu_pa_msg[21]),
	.msg_out_22      (cnu_pa_msg[22]),
	.msg_out_23      (cnu_pa_msg[23]),
	.msg_out_24      (cnu_pa_msg[24]),
	.msg_out_25      (cnu_pa_msg[25]),
	.msg_out_26      (cnu_pa_msg[26]),
	.msg_out_27      (cnu_pa_msg[27]),
	.msg_out_28      (cnu_pa_msg[28]),
	.msg_out_29      (cnu_pa_msg[29]),
	.msg_out_30      (cnu_pa_msg[30]),
	.msg_out_31      (cnu_pa_msg[31]),
	.msg_out_32      (cnu_pa_msg[32]),
	.msg_out_33      (cnu_pa_msg[33]),
	.msg_out_34      (cnu_pa_msg[34]),
	.msg_out_35      (cnu_pa_msg[35]),
	.msg_out_36      (cnu_pa_msg[36]),
	.msg_out_37      (cnu_pa_msg[37]),
	.msg_out_38      (cnu_pa_msg[38]),
	.msg_out_39      (cnu_pa_msg[39]),
	.msg_out_40      (cnu_pa_msg[40]),
	.msg_out_41      (cnu_pa_msg[41]),
	.msg_out_42      (cnu_pa_msg[42]),
	.msg_out_43      (cnu_pa_msg[43]),
	.msg_out_44      (cnu_pa_msg[44]),
	.msg_out_45      (cnu_pa_msg[45]),
	.msg_out_46      (cnu_pa_msg[46]),
	.msg_out_47      (cnu_pa_msg[47]),
	.msg_out_48      (cnu_pa_msg[48]),
	.msg_out_49      (cnu_pa_msg[49]),
	.msg_out_50      (cnu_pa_msg[50]),
	.msg_out_51      (cnu_pa_msg[51]),
	.msg_out_52      (cnu_pa_msg[52]),
	.msg_out_53      (cnu_pa_msg[53]),
	.msg_out_54      (cnu_pa_msg[54]),
	.msg_out_55      (cnu_pa_msg[55]),
	.msg_out_56      (cnu_pa_msg[56]),
	.msg_out_57      (cnu_pa_msg[57]),
	.msg_out_58      (cnu_pa_msg[58]),
	.msg_out_59      (cnu_pa_msg[59]),
	.msg_out_60      (cnu_pa_msg[60]),
	.msg_out_61      (cnu_pa_msg[61]),
	.msg_out_62      (cnu_pa_msg[62]),
	.msg_out_63      (cnu_pa_msg[63]),
	.msg_out_64      (cnu_pa_msg[64]),
	.msg_out_65      (cnu_pa_msg[65]),
	.msg_out_66      (cnu_pa_msg[66]),
	.msg_out_67      (cnu_pa_msg[67]),
	.msg_out_68      (cnu_pa_msg[68]),
	.msg_out_69      (cnu_pa_msg[69]),
	.msg_out_70      (cnu_pa_msg[70]),
	.msg_out_71      (cnu_pa_msg[71]),
	.msg_out_72      (cnu_pa_msg[72]),
	.msg_out_73      (cnu_pa_msg[73]),
	.msg_out_74      (cnu_pa_msg[74]),
	.msg_out_75      (cnu_pa_msg[75]),
	.msg_out_76      (cnu_pa_msg[76]),
	.msg_out_77      (cnu_pa_msg[77]),
	.msg_out_78      (cnu_pa_msg[78]),
	.msg_out_79      (cnu_pa_msg[79]),
	.msg_out_80      (cnu_pa_msg[80]),
	.msg_out_81      (cnu_pa_msg[81]),
	.msg_out_82      (cnu_pa_msg[82]),
	.msg_out_83      (cnu_pa_msg[83]),
	.msg_out_84      (cnu_pa_msg[84]),
	.msg_in_0        (cnu_to_mem_0),
	.msg_in_1        (cnu_to_mem_1),
	.msg_in_2        (cnu_to_mem_2),
	.msg_in_3        (cnu_to_mem_3),
	.msg_in_4        (cnu_to_mem_4),
	.msg_in_5        (cnu_to_mem_5),
	.msg_in_6        (cnu_to_mem_6),
	.msg_in_7        (cnu_to_mem_7),
	.msg_in_8        (cnu_to_mem_8),
	.msg_in_9        (cnu_to_mem_9),
	.msg_in_10       (cnu_to_mem_10),
	.msg_in_11       (cnu_to_mem_11),
	.msg_in_12       (cnu_to_mem_12),
	.msg_in_13       (cnu_to_mem_13),
	.msg_in_14       (cnu_to_mem_14),
	.msg_in_15       (cnu_to_mem_15),
	.msg_in_16       (cnu_to_mem_16),
	.msg_in_17       (cnu_to_mem_17),
	.msg_in_18       (cnu_to_mem_18),
	.msg_in_19       (cnu_to_mem_19),
	.msg_in_20       (cnu_to_mem_20),
	.msg_in_21       (cnu_to_mem_21),
	.msg_in_22       (cnu_to_mem_22),
	.msg_in_23       (cnu_to_mem_23),
	.msg_in_24       (cnu_to_mem_24),
	.msg_in_25       (cnu_to_mem_25),
	.msg_in_26       (cnu_to_mem_26),
	.msg_in_27       (cnu_to_mem_27),
	.msg_in_28       (cnu_to_mem_28),
	.msg_in_29       (cnu_to_mem_29),
	.msg_in_30       (cnu_to_mem_30),
	.msg_in_31       (cnu_to_mem_31),
	.msg_in_32       (cnu_to_mem_32),
	.msg_in_33       (cnu_to_mem_33),
	.msg_in_34       (cnu_to_mem_34),
	.msg_in_35       (cnu_to_mem_35),
	.msg_in_36       (cnu_to_mem_36),
	.msg_in_37       (cnu_to_mem_37),
	.msg_in_38       (cnu_to_mem_38),
	.msg_in_39       (cnu_to_mem_39),
	.msg_in_40       (cnu_to_mem_40),
	.msg_in_41       (cnu_to_mem_41),
	.msg_in_42       (cnu_to_mem_42),
	.msg_in_43       (cnu_to_mem_43),
	.msg_in_44       (cnu_to_mem_44),
	.msg_in_45       (cnu_to_mem_45),
	.msg_in_46       (cnu_to_mem_46),
	.msg_in_47       (cnu_to_mem_47),
	.msg_in_48       (cnu_to_mem_48),
	.msg_in_49       (cnu_to_mem_49),
	.msg_in_50       (cnu_to_mem_50),
	.msg_in_51       (cnu_to_mem_51),
	.msg_in_52       (cnu_to_mem_52),
	.msg_in_53       (cnu_to_mem_53),
	.msg_in_54       (cnu_to_mem_54),
	.msg_in_55       (cnu_to_mem_55),
	.msg_in_56       (cnu_to_mem_56),
	.msg_in_57       (cnu_to_mem_57),
	.msg_in_58       (cnu_to_mem_58),
	.msg_in_59       (cnu_to_mem_59),
	.msg_in_60       (cnu_to_mem_60),
	.msg_in_61       (cnu_to_mem_61),
	.msg_in_62       (cnu_to_mem_62),
	.msg_in_63       (cnu_to_mem_63),
	.msg_in_64       (cnu_to_mem_64),
	.msg_in_65       (cnu_to_mem_65),
	.msg_in_66       (cnu_to_mem_66),
	.msg_in_67       (cnu_to_mem_67),
	.msg_in_68       (cnu_to_mem_68),
	.msg_in_69       (cnu_to_mem_69),
	.msg_in_70       (cnu_to_mem_70),
	.msg_in_71       (cnu_to_mem_71),
	.msg_in_72       (cnu_to_mem_72),
	.msg_in_73       (cnu_to_mem_73),
	.msg_in_74       (cnu_to_mem_74),
	.msg_in_75       (cnu_to_mem_75),
	.msg_in_76       (cnu_to_mem_76),
	.msg_in_77       (cnu_to_mem_77),
	.msg_in_78       (cnu_to_mem_78),
	.msg_in_79       (cnu_to_mem_79),
	.msg_in_80       (cnu_to_mem_80),
	.msg_in_81       (cnu_to_mem_81),
	.msg_in_82       (cnu_to_mem_82),
	.msg_in_83       (cnu_to_mem_83),
	.msg_in_84       (cnu_to_mem_84),
	.layer_status    (cnu_layer_status),
	.first_row_chunk (last_row_chunk[0]),
	.sys_clk         (sys_clk),
	.rstn            (rstn)
);
/*-------------------------------------------------------*/
// Page alignment of Variable nodes
wire [QUAN_SIZE-1:0] vnu_pa_msg [CHECK_PARALLELISM-1:0];
ram_pageAlign_interface_submatrix_9 #(
	.QUAN_SIZE(QUAN_SIZE),
	.CHECK_PARALLELISM(CHECK_PARALLELISM),
	.LAYER_NUM(LAYER_NUM)
) vnu_ram_pageAlign_interface_submatrix_9 (
	.msg_out_0       (vnu_pa_msg[0 ]),
	.msg_out_1       (vnu_pa_msg[1 ]),
	.msg_out_2       (vnu_pa_msg[2 ]),
	.msg_out_3       (vnu_pa_msg[3 ]),
	.msg_out_4       (vnu_pa_msg[4 ]),
	.msg_out_5       (vnu_pa_msg[5 ]),
	.msg_out_6       (vnu_pa_msg[6 ]),
	.msg_out_7       (vnu_pa_msg[7 ]),
	.msg_out_8       (vnu_pa_msg[8 ]),
	.msg_out_9       (vnu_pa_msg[9 ]),
	.msg_out_10      (vnu_pa_msg[10]),
	.msg_out_11      (vnu_pa_msg[11]),
	.msg_out_12      (vnu_pa_msg[12]),
	.msg_out_13      (vnu_pa_msg[13]),
	.msg_out_14      (vnu_pa_msg[14]),
	.msg_out_15      (vnu_pa_msg[15]),
	.msg_out_16      (vnu_pa_msg[16]),
	.msg_out_17      (vnu_pa_msg[17]),
	.msg_out_18      (vnu_pa_msg[18]),
	.msg_out_19      (vnu_pa_msg[19]),
	.msg_out_20      (vnu_pa_msg[20]),
	.msg_out_21      (vnu_pa_msg[21]),
	.msg_out_22      (vnu_pa_msg[22]),
	.msg_out_23      (vnu_pa_msg[23]),
	.msg_out_24      (vnu_pa_msg[24]),
	.msg_out_25      (vnu_pa_msg[25]),
	.msg_out_26      (vnu_pa_msg[26]),
	.msg_out_27      (vnu_pa_msg[27]),
	.msg_out_28      (vnu_pa_msg[28]),
	.msg_out_29      (vnu_pa_msg[29]),
	.msg_out_30      (vnu_pa_msg[30]),
	.msg_out_31      (vnu_pa_msg[31]),
	.msg_out_32      (vnu_pa_msg[32]),
	.msg_out_33      (vnu_pa_msg[33]),
	.msg_out_34      (vnu_pa_msg[34]),
	.msg_out_35      (vnu_pa_msg[35]),
	.msg_out_36      (vnu_pa_msg[36]),
	.msg_out_37      (vnu_pa_msg[37]),
	.msg_out_38      (vnu_pa_msg[38]),
	.msg_out_39      (vnu_pa_msg[39]),
	.msg_out_40      (vnu_pa_msg[40]),
	.msg_out_41      (vnu_pa_msg[41]),
	.msg_out_42      (vnu_pa_msg[42]),
	.msg_out_43      (vnu_pa_msg[43]),
	.msg_out_44      (vnu_pa_msg[44]),
	.msg_out_45      (vnu_pa_msg[45]),
	.msg_out_46      (vnu_pa_msg[46]),
	.msg_out_47      (vnu_pa_msg[47]),
	.msg_out_48      (vnu_pa_msg[48]),
	.msg_out_49      (vnu_pa_msg[49]),
	.msg_out_50      (vnu_pa_msg[50]),
	.msg_out_51      (vnu_pa_msg[51]),
	.msg_out_52      (vnu_pa_msg[52]),
	.msg_out_53      (vnu_pa_msg[53]),
	.msg_out_54      (vnu_pa_msg[54]),
	.msg_out_55      (vnu_pa_msg[55]),
	.msg_out_56      (vnu_pa_msg[56]),
	.msg_out_57      (vnu_pa_msg[57]),
	.msg_out_58      (vnu_pa_msg[58]),
	.msg_out_59      (vnu_pa_msg[59]),
	.msg_out_60      (vnu_pa_msg[60]),
	.msg_out_61      (vnu_pa_msg[61]),
	.msg_out_62      (vnu_pa_msg[62]),
	.msg_out_63      (vnu_pa_msg[63]),
	.msg_out_64      (vnu_pa_msg[64]),
	.msg_out_65      (vnu_pa_msg[65]),
	.msg_out_66      (vnu_pa_msg[66]),
	.msg_out_67      (vnu_pa_msg[67]),
	.msg_out_68      (vnu_pa_msg[68]),
	.msg_out_69      (vnu_pa_msg[69]),
	.msg_out_70      (vnu_pa_msg[70]),
	.msg_out_71      (vnu_pa_msg[71]),
	.msg_out_72      (vnu_pa_msg[72]),
	.msg_out_73      (vnu_pa_msg[73]),
	.msg_out_74      (vnu_pa_msg[74]),
	.msg_out_75      (vnu_pa_msg[75]),
	.msg_out_76      (vnu_pa_msg[76]),
	.msg_out_77      (vnu_pa_msg[77]),
	.msg_out_78      (vnu_pa_msg[78]),
	.msg_out_79      (vnu_pa_msg[79]),
	.msg_out_80      (vnu_pa_msg[80]),
	.msg_out_81      (vnu_pa_msg[81]),
	.msg_out_82      (vnu_pa_msg[82]),
	.msg_out_83      (vnu_pa_msg[83]),
	.msg_out_84      (vnu_pa_msg[84]),
	.msg_in_0        (vnu_to_mem_0),
	.msg_in_1        (vnu_to_mem_1),
	.msg_in_2        (vnu_to_mem_2),
	.msg_in_3        (vnu_to_mem_3),
	.msg_in_4        (vnu_to_mem_4),
	.msg_in_5        (vnu_to_mem_5),
	.msg_in_6        (vnu_to_mem_6),
	.msg_in_7        (vnu_to_mem_7),
	.msg_in_8        (vnu_to_mem_8),
	.msg_in_9        (vnu_to_mem_9),
	.msg_in_10       (vnu_to_mem_10),
	.msg_in_11       (vnu_to_mem_11),
	.msg_in_12       (vnu_to_mem_12),
	.msg_in_13       (vnu_to_mem_13),
	.msg_in_14       (vnu_to_mem_14),
	.msg_in_15       (vnu_to_mem_15),
	.msg_in_16       (vnu_to_mem_16),
	.msg_in_17       (vnu_to_mem_17),
	.msg_in_18       (vnu_to_mem_18),
	.msg_in_19       (vnu_to_mem_19),
	.msg_in_20       (vnu_to_mem_20),
	.msg_in_21       (vnu_to_mem_21),
	.msg_in_22       (vnu_to_mem_22),
	.msg_in_23       (vnu_to_mem_23),
	.msg_in_24       (vnu_to_mem_24),
	.msg_in_25       (vnu_to_mem_25),
	.msg_in_26       (vnu_to_mem_26),
	.msg_in_27       (vnu_to_mem_27),
	.msg_in_28       (vnu_to_mem_28),
	.msg_in_29       (vnu_to_mem_29),
	.msg_in_30       (vnu_to_mem_30),
	.msg_in_31       (vnu_to_mem_31),
	.msg_in_32       (vnu_to_mem_32),
	.msg_in_33       (vnu_to_mem_33),
	.msg_in_34       (vnu_to_mem_34),
	.msg_in_35       (vnu_to_mem_35),
	.msg_in_36       (vnu_to_mem_36),
	.msg_in_37       (vnu_to_mem_37),
	.msg_in_38       (vnu_to_mem_38),
	.msg_in_39       (vnu_to_mem_39),
	.msg_in_40       (vnu_to_mem_40),
	.msg_in_41       (vnu_to_mem_41),
	.msg_in_42       (vnu_to_mem_42),
	.msg_in_43       (vnu_to_mem_43),
	.msg_in_44       (vnu_to_mem_44),
	.msg_in_45       (vnu_to_mem_45),
	.msg_in_46       (vnu_to_mem_46),
	.msg_in_47       (vnu_to_mem_47),
	.msg_in_48       (vnu_to_mem_48),
	.msg_in_49       (vnu_to_mem_49),
	.msg_in_50       (vnu_to_mem_50),
	.msg_in_51       (vnu_to_mem_51),
	.msg_in_52       (vnu_to_mem_52),
	.msg_in_53       (vnu_to_mem_53),
	.msg_in_54       (vnu_to_mem_54),
	.msg_in_55       (vnu_to_mem_55),
	.msg_in_56       (vnu_to_mem_56),
	.msg_in_57       (vnu_to_mem_57),
	.msg_in_58       (vnu_to_mem_58),
	.msg_in_59       (vnu_to_mem_59),
	.msg_in_60       (vnu_to_mem_60),
	.msg_in_61       (vnu_to_mem_61),
	.msg_in_62       (vnu_to_mem_62),
	.msg_in_63       (vnu_to_mem_63),
	.msg_in_64       (vnu_to_mem_64),
	.msg_in_65       (vnu_to_mem_65),
	.msg_in_66       (vnu_to_mem_66),
	.msg_in_67       (vnu_to_mem_67),
	.msg_in_68       (vnu_to_mem_68),
	.msg_in_69       (vnu_to_mem_69),
	.msg_in_70       (vnu_to_mem_70),
	.msg_in_71       (vnu_to_mem_71),
	.msg_in_72       (vnu_to_mem_72),
	.msg_in_73       (vnu_to_mem_73),
	.msg_in_74       (vnu_to_mem_74),
	.msg_in_75       (vnu_to_mem_75),
	.msg_in_76       (vnu_to_mem_76),
	.msg_in_77       (vnu_to_mem_77),
	.msg_in_78       (vnu_to_mem_78),
	.msg_in_79       (vnu_to_mem_79),
	.msg_in_80       (vnu_to_mem_80),
	.msg_in_81       (vnu_to_mem_81),
	.msg_in_82       (vnu_to_mem_82),
	.msg_in_83       (vnu_to_mem_83),
	.msg_in_84       (vnu_to_mem_84),
	.layer_status    (vnu_layer_status),
	.first_row_chunk (last_row_chunk[1]),
	.sys_clk         (sys_clk),
	.rstn            (rstn)
);
/*-------------------------------------------------------*/
// Memory Instantiation
column_ram_pc85 #(
	.QUAN_SIZE(QUAN_SIZE),
	.CHECK_PARALLELISM(CHECK_PARALLELISM),
	.RAM_PORTA_RANGE(RAM_PORTA_RANGE),
	.RAM_PORTB_RANGE(RAM_PORTB_RANGE),
	.MEM_DEVICE_NUM(MEM_DEVICE_NUM),
	.DEPTH(DEPTH),
	.DATA_WIDTH(DATA_WIDTH),
	.FRAG_DATA_WIDTH(FRAG_DATA_WIDTH),
	.ADDR_WIDTH(ADDR_WIDTH)
) inst_column_ram_pc85 (
	.first_dout_0   (mem_to_cnu_0 ),
	.first_dout_1   (mem_to_cnu_1 ),
	.first_dout_2   (mem_to_cnu_2 ),
	.first_dout_3   (mem_to_cnu_3 ),
	.first_dout_4   (mem_to_cnu_4 ),
	.first_dout_5   (mem_to_cnu_5 ),
	.first_dout_6   (mem_to_cnu_6 ),
	.first_dout_7   (mem_to_cnu_7 ),
	.first_dout_8   (mem_to_cnu_8 ),
	.first_dout_9   (mem_to_cnu_9 ),
	.first_dout_10  (mem_to_cnu_10),
	.first_dout_11  (mem_to_cnu_11),
	.first_dout_12  (mem_to_cnu_12),
	.first_dout_13  (mem_to_cnu_13),
	.first_dout_14  (mem_to_cnu_14),
	.first_dout_15  (mem_to_cnu_15),
	.first_dout_16  (mem_to_cnu_16),
	.first_dout_17  (mem_to_cnu_17),
	.first_dout_18  (mem_to_cnu_18),
	.first_dout_19  (mem_to_cnu_19),
	.first_dout_20  (mem_to_cnu_20),
	.first_dout_21  (mem_to_cnu_21),
	.first_dout_22  (mem_to_cnu_22),
	.first_dout_23  (mem_to_cnu_23),
	.first_dout_24  (mem_to_cnu_24),
	.first_dout_25  (mem_to_cnu_25),
	.first_dout_26  (mem_to_cnu_26),
	.first_dout_27  (mem_to_cnu_27),
	.first_dout_28  (mem_to_cnu_28),
	.first_dout_29  (mem_to_cnu_29),
	.first_dout_30  (mem_to_cnu_30),
	.first_dout_31  (mem_to_cnu_31),
	.first_dout_32  (mem_to_cnu_32),
	.first_dout_33  (mem_to_cnu_33),
	.first_dout_34  (mem_to_cnu_34),
	.first_dout_35  (mem_to_cnu_35),
	.first_dout_36  (mem_to_cnu_36),
	.first_dout_37  (mem_to_cnu_37),
	.first_dout_38  (mem_to_cnu_38),
	.first_dout_39  (mem_to_cnu_39),
	.first_dout_40  (mem_to_cnu_40),
	.first_dout_41  (mem_to_cnu_41),
	.first_dout_42  (mem_to_cnu_42),
	.first_dout_43  (mem_to_cnu_43),
	.first_dout_44  (mem_to_cnu_44),
	.first_dout_45  (mem_to_cnu_45),
	.first_dout_46  (mem_to_cnu_46),
	.first_dout_47  (mem_to_cnu_47),
	.first_dout_48  (mem_to_cnu_48),
	.first_dout_49  (mem_to_cnu_49),
	.first_dout_50  (mem_to_cnu_50),
	.first_dout_51  (mem_to_cnu_51),
	.first_dout_52  (mem_to_cnu_52),
	.first_dout_53  (mem_to_cnu_53),
	.first_dout_54  (mem_to_cnu_54),
	.first_dout_55  (mem_to_cnu_55),
	.first_dout_56  (mem_to_cnu_56),
	.first_dout_57  (mem_to_cnu_57),
	.first_dout_58  (mem_to_cnu_58),
	.first_dout_59  (mem_to_cnu_59),
	.first_dout_60  (mem_to_cnu_60),
	.first_dout_61  (mem_to_cnu_61),
	.first_dout_62  (mem_to_cnu_62),
	.first_dout_63  (mem_to_cnu_63),
	.first_dout_64  (mem_to_cnu_64),
	.first_dout_65  (mem_to_cnu_65),
	.first_dout_66  (mem_to_cnu_66),
	.first_dout_67  (mem_to_cnu_67),
	.first_dout_68  (mem_to_cnu_68),
	.first_dout_69  (mem_to_cnu_69),
	.first_dout_70  (mem_to_cnu_70),
	.first_dout_71  (mem_to_cnu_71),
	.first_dout_72  (mem_to_cnu_72),
	.first_dout_73  (mem_to_cnu_73),
	.first_dout_74  (mem_to_cnu_74),
	.first_dout_75  (mem_to_cnu_75),
	.first_dout_76  (mem_to_cnu_76),
	.first_dout_77  (mem_to_cnu_77),
	.first_dout_78  (mem_to_cnu_78),
	.first_dout_79  (mem_to_cnu_79),
	.first_dout_80  (mem_to_cnu_80),
	.first_dout_81  (mem_to_cnu_81),
	.first_dout_82  (mem_to_cnu_82),
	.first_dout_83  (mem_to_cnu_83),
	.first_dout_84  (mem_to_cnu_84),
	.second_dout_0  (mem_to_vnu_0 ),
	.second_dout_1  (mem_to_vnu_1 ),
	.second_dout_2  (mem_to_vnu_2 ),
	.second_dout_3  (mem_to_vnu_3 ),
	.second_dout_4  (mem_to_vnu_4 ),
	.second_dout_5  (mem_to_vnu_5 ),
	.second_dout_6  (mem_to_vnu_6 ),
	.second_dout_7  (mem_to_vnu_7 ),
	.second_dout_8  (mem_to_vnu_8 ),
	.second_dout_9  (mem_to_vnu_9 ),
	.second_dout_10 (mem_to_vnu_10),
	.second_dout_11 (mem_to_vnu_11),
	.second_dout_12 (mem_to_vnu_12),
	.second_dout_13 (mem_to_vnu_13),
	.second_dout_14 (mem_to_vnu_14),
	.second_dout_15 (mem_to_vnu_15),
	.second_dout_16 (mem_to_vnu_16),
	.second_dout_17 (mem_to_vnu_17),
	.second_dout_18 (mem_to_vnu_18),
	.second_dout_19 (mem_to_vnu_19),
	.second_dout_20 (mem_to_vnu_20),
	.second_dout_21 (mem_to_vnu_21),
	.second_dout_22 (mem_to_vnu_22),
	.second_dout_23 (mem_to_vnu_23),
	.second_dout_24 (mem_to_vnu_24),
	.second_dout_25 (mem_to_vnu_25),
	.second_dout_26 (mem_to_vnu_26),
	.second_dout_27 (mem_to_vnu_27),
	.second_dout_28 (mem_to_vnu_28),
	.second_dout_29 (mem_to_vnu_29),
	.second_dout_30 (mem_to_vnu_30),
	.second_dout_31 (mem_to_vnu_31),
	.second_dout_32 (mem_to_vnu_32),
	.second_dout_33 (mem_to_vnu_33),
	.second_dout_34 (mem_to_vnu_34),
	.second_dout_35 (mem_to_vnu_35),
	.second_dout_36 (mem_to_vnu_36),
	.second_dout_37 (mem_to_vnu_37),
	.second_dout_38 (mem_to_vnu_38),
	.second_dout_39 (mem_to_vnu_39),
	.second_dout_40 (mem_to_vnu_40),
	.second_dout_41 (mem_to_vnu_41),
	.second_dout_42 (mem_to_vnu_42),
	.second_dout_43 (mem_to_vnu_43),
	.second_dout_44 (mem_to_vnu_44),
	.second_dout_45 (mem_to_vnu_45),
	.second_dout_46 (mem_to_vnu_46),
	.second_dout_47 (mem_to_vnu_47),
	.second_dout_48 (mem_to_vnu_48),
	.second_dout_49 (mem_to_vnu_49),
	.second_dout_50 (mem_to_vnu_50),
	.second_dout_51 (mem_to_vnu_51),
	.second_dout_52 (mem_to_vnu_52),
	.second_dout_53 (mem_to_vnu_53),
	.second_dout_54 (mem_to_vnu_54),
	.second_dout_55 (mem_to_vnu_55),
	.second_dout_56 (mem_to_vnu_56),
	.second_dout_57 (mem_to_vnu_57),
	.second_dout_58 (mem_to_vnu_58),
	.second_dout_59 (mem_to_vnu_59),
	.second_dout_60 (mem_to_vnu_60),
	.second_dout_61 (mem_to_vnu_61),
	.second_dout_62 (mem_to_vnu_62),
	.second_dout_63 (mem_to_vnu_63),
	.second_dout_64 (mem_to_vnu_64),
	.second_dout_65 (mem_to_vnu_65),
	.second_dout_66 (mem_to_vnu_66),
	.second_dout_67 (mem_to_vnu_67),
	.second_dout_68 (mem_to_vnu_68),
	.second_dout_69 (mem_to_vnu_69),
	.second_dout_70 (mem_to_vnu_70),
	.second_dout_71 (mem_to_vnu_71),
	.second_dout_72 (mem_to_vnu_72),
	.second_dout_73 (mem_to_vnu_73),
	.second_dout_74 (mem_to_vnu_74),
	.second_dout_75 (mem_to_vnu_75),
	.second_dout_76 (mem_to_vnu_76),
	.second_dout_77 (mem_to_vnu_77),
	.second_dout_78 (mem_to_vnu_78),
	.second_dout_79 (mem_to_vnu_79),
	.second_dout_80 (mem_to_vnu_80),
	.second_dout_81 (mem_to_vnu_81),
	.second_dout_82 (mem_to_vnu_82),
	.second_dout_83 (mem_to_vnu_83),
	.second_dout_84 (mem_to_vnu_84),
	.first_din_0    (cnu_pa_msg[0 ]),
	.first_din_1    (cnu_pa_msg[1 ]),
	.first_din_2    (cnu_pa_msg[2 ]),
	.first_din_3    (cnu_pa_msg[3 ]),
	.first_din_4    (cnu_pa_msg[4 ]),
	.first_din_5    (cnu_pa_msg[5 ]),
	.first_din_6    (cnu_pa_msg[6 ]),
	.first_din_7    (cnu_pa_msg[7 ]),
	.first_din_8    (cnu_pa_msg[8 ]),
	.first_din_9    (cnu_pa_msg[9 ]),
	.first_din_10   (cnu_pa_msg[10]),
	.first_din_11   (cnu_pa_msg[11]),
	.first_din_12   (cnu_pa_msg[12]),
	.first_din_13   (cnu_pa_msg[13]),
	.first_din_14   (cnu_pa_msg[14]),
	.first_din_15   (cnu_pa_msg[15]),
	.first_din_16   (cnu_pa_msg[16]),
	.first_din_17   (cnu_pa_msg[17]),
	.first_din_18   (cnu_pa_msg[18]),
	.first_din_19   (cnu_pa_msg[19]),
	.first_din_20   (cnu_pa_msg[20]),
	.first_din_21   (cnu_pa_msg[21]),
	.first_din_22   (cnu_pa_msg[22]),
	.first_din_23   (cnu_pa_msg[23]),
	.first_din_24   (cnu_pa_msg[24]),
	.first_din_25   (cnu_pa_msg[25]),
	.first_din_26   (cnu_pa_msg[26]),
	.first_din_27   (cnu_pa_msg[27]),
	.first_din_28   (cnu_pa_msg[28]),
	.first_din_29   (cnu_pa_msg[29]),
	.first_din_30   (cnu_pa_msg[30]),
	.first_din_31   (cnu_pa_msg[31]),
	.first_din_32   (cnu_pa_msg[32]),
	.first_din_33   (cnu_pa_msg[33]),
	.first_din_34   (cnu_pa_msg[34]),
	.first_din_35   (cnu_pa_msg[35]),
	.first_din_36   (cnu_pa_msg[36]),
	.first_din_37   (cnu_pa_msg[37]),
	.first_din_38   (cnu_pa_msg[38]),
	.first_din_39   (cnu_pa_msg[39]),
	.first_din_40   (cnu_pa_msg[40]),
	.first_din_41   (cnu_pa_msg[41]),
	.first_din_42   (cnu_pa_msg[42]),
	.first_din_43   (cnu_pa_msg[43]),
	.first_din_44   (cnu_pa_msg[44]),
	.first_din_45   (cnu_pa_msg[45]),
	.first_din_46   (cnu_pa_msg[46]),
	.first_din_47   (cnu_pa_msg[47]),
	.first_din_48   (cnu_pa_msg[48]),
	.first_din_49   (cnu_pa_msg[49]),
	.first_din_50   (cnu_pa_msg[50]),
	.first_din_51   (cnu_pa_msg[51]),
	.first_din_52   (cnu_pa_msg[52]),
	.first_din_53   (cnu_pa_msg[53]),
	.first_din_54   (cnu_pa_msg[54]),
	.first_din_55   (cnu_pa_msg[55]),
	.first_din_56   (cnu_pa_msg[56]),
	.first_din_57   (cnu_pa_msg[57]),
	.first_din_58   (cnu_pa_msg[58]),
	.first_din_59   (cnu_pa_msg[59]),
	.first_din_60   (cnu_pa_msg[60]),
	.first_din_61   (cnu_pa_msg[61]),
	.first_din_62   (cnu_pa_msg[62]),
	.first_din_63   (cnu_pa_msg[63]),
	.first_din_64   (cnu_pa_msg[64]),
	.first_din_65   (cnu_pa_msg[65]),
	.first_din_66   (cnu_pa_msg[66]),
	.first_din_67   (cnu_pa_msg[67]),
	.first_din_68   (cnu_pa_msg[68]),
	.first_din_69   (cnu_pa_msg[69]),
	.first_din_70   (cnu_pa_msg[70]),
	.first_din_71   (cnu_pa_msg[71]),
	.first_din_72   (cnu_pa_msg[72]),
	.first_din_73   (cnu_pa_msg[73]),
	.first_din_74   (cnu_pa_msg[74]),
	.first_din_75   (cnu_pa_msg[75]),
	.first_din_76   (cnu_pa_msg[76]),
	.first_din_77   (cnu_pa_msg[77]),
	.first_din_78   (cnu_pa_msg[78]),
	.first_din_79   (cnu_pa_msg[79]),
	.first_din_80   (cnu_pa_msg[80]),
	.first_din_81   (cnu_pa_msg[81]),
	.first_din_82   (cnu_pa_msg[82]),
	.first_din_83   (cnu_pa_msg[83]),
	.first_din_84   (cnu_pa_msg[84]),
	.second_din_0   (vnu_pa_msg[0 ]),
	.second_din_1   (vnu_pa_msg[1 ]),
	.second_din_2   (vnu_pa_msg[2 ]),
	.second_din_3   (vnu_pa_msg[3 ]),
	.second_din_4   (vnu_pa_msg[4 ]),
	.second_din_5   (vnu_pa_msg[5 ]),
	.second_din_6   (vnu_pa_msg[6 ]),
	.second_din_7   (vnu_pa_msg[7 ]),
	.second_din_8   (vnu_pa_msg[8 ]),
	.second_din_9   (vnu_pa_msg[9 ]),
	.second_din_10  (vnu_pa_msg[10]),
	.second_din_11  (vnu_pa_msg[11]),
	.second_din_12  (vnu_pa_msg[12]),
	.second_din_13  (vnu_pa_msg[13]),
	.second_din_14  (vnu_pa_msg[14]),
	.second_din_15  (vnu_pa_msg[15]),
	.second_din_16  (vnu_pa_msg[16]),
	.second_din_17  (vnu_pa_msg[17]),
	.second_din_18  (vnu_pa_msg[18]),
	.second_din_19  (vnu_pa_msg[19]),
	.second_din_20  (vnu_pa_msg[20]),
	.second_din_21  (vnu_pa_msg[21]),
	.second_din_22  (vnu_pa_msg[22]),
	.second_din_23  (vnu_pa_msg[23]),
	.second_din_24  (vnu_pa_msg[24]),
	.second_din_25  (vnu_pa_msg[25]),
	.second_din_26  (vnu_pa_msg[26]),
	.second_din_27  (vnu_pa_msg[27]),
	.second_din_28  (vnu_pa_msg[28]),
	.second_din_29  (vnu_pa_msg[29]),
	.second_din_30  (vnu_pa_msg[30]),
	.second_din_31  (vnu_pa_msg[31]),
	.second_din_32  (vnu_pa_msg[32]),
	.second_din_33  (vnu_pa_msg[33]),
	.second_din_34  (vnu_pa_msg[34]),
	.second_din_35  (vnu_pa_msg[35]),
	.second_din_36  (vnu_pa_msg[36]),
	.second_din_37  (vnu_pa_msg[37]),
	.second_din_38  (vnu_pa_msg[38]),
	.second_din_39  (vnu_pa_msg[39]),
	.second_din_40  (vnu_pa_msg[40]),
	.second_din_41  (vnu_pa_msg[41]),
	.second_din_42  (vnu_pa_msg[42]),
	.second_din_43  (vnu_pa_msg[43]),
	.second_din_44  (vnu_pa_msg[44]),
	.second_din_45  (vnu_pa_msg[45]),
	.second_din_46  (vnu_pa_msg[46]),
	.second_din_47  (vnu_pa_msg[47]),
	.second_din_48  (vnu_pa_msg[48]),
	.second_din_49  (vnu_pa_msg[49]),
	.second_din_50  (vnu_pa_msg[50]),
	.second_din_51  (vnu_pa_msg[51]),
	.second_din_52  (vnu_pa_msg[52]),
	.second_din_53  (vnu_pa_msg[53]),
	.second_din_54  (vnu_pa_msg[54]),
	.second_din_55  (vnu_pa_msg[55]),
	.second_din_56  (vnu_pa_msg[56]),
	.second_din_57  (vnu_pa_msg[57]),
	.second_din_58  (vnu_pa_msg[58]),
	.second_din_59  (vnu_pa_msg[59]),
	.second_din_60  (vnu_pa_msg[60]),
	.second_din_61  (vnu_pa_msg[61]),
	.second_din_62  (vnu_pa_msg[62]),
	.second_din_63  (vnu_pa_msg[63]),
	.second_din_64  (vnu_pa_msg[64]),
	.second_din_65  (vnu_pa_msg[65]),
	.second_din_66  (vnu_pa_msg[66]),
	.second_din_67  (vnu_pa_msg[67]),
	.second_din_68  (vnu_pa_msg[68]),
	.second_din_69  (vnu_pa_msg[69]),
	.second_din_70  (vnu_pa_msg[70]),
	.second_din_71  (vnu_pa_msg[71]),
	.second_din_72  (vnu_pa_msg[72]),
	.second_din_73  (vnu_pa_msg[73]),
	.second_din_74  (vnu_pa_msg[74]),
	.second_din_75  (vnu_pa_msg[75]),
	.second_din_76  (vnu_pa_msg[76]),
	.second_din_77  (vnu_pa_msg[77]),
	.second_din_78  (vnu_pa_msg[78]),
	.second_din_79  (vnu_pa_msg[79]),
	.second_din_80  (vnu_pa_msg[80]),
	.second_din_81  (vnu_pa_msg[81]),
	.second_din_82  (vnu_pa_msg[82]),
	.second_din_83  (vnu_pa_msg[83]),
	.second_din_84  (vnu_pa_msg[84]),

	.sync_addr_0    (cnu_sync_addr),
	.sync_addr_1    (vnu_sync_addr),
	.we             (we),
	.sys_clk        (sys_clk)
);
assign vnu_pa_msg_bit0[CHECK_PARALLELISM-1:0] = {vnu_pa_msg[84][0],vnu_pa_msg[83][0],vnu_pa_msg[82][0],vnu_pa_msg[81][0],vnu_pa_msg[80][0],vnu_pa_msg[79][0],vnu_pa_msg[78][0],vnu_pa_msg[77][0],vnu_pa_msg[76][0],vnu_pa_msg[75][0],vnu_pa_msg[74][0],vnu_pa_msg[73][0],vnu_pa_msg[72][0],vnu_pa_msg[71][0],vnu_pa_msg[70][0],vnu_pa_msg[69][0],vnu_pa_msg[68][0],vnu_pa_msg[67][0],vnu_pa_msg[66][0],vnu_pa_msg[65][0],vnu_pa_msg[64][0],vnu_pa_msg[63][0],vnu_pa_msg[62][0],vnu_pa_msg[61][0],vnu_pa_msg[60][0],vnu_pa_msg[59][0],vnu_pa_msg[58][0],vnu_pa_msg[57][0],vnu_pa_msg[56][0],vnu_pa_msg[55][0],vnu_pa_msg[54][0],vnu_pa_msg[53][0],vnu_pa_msg[52][0],vnu_pa_msg[51][0],vnu_pa_msg[50][0],vnu_pa_msg[49][0],vnu_pa_msg[48][0],vnu_pa_msg[47][0],vnu_pa_msg[46][0],vnu_pa_msg[45][0],vnu_pa_msg[44][0],vnu_pa_msg[43][0],vnu_pa_msg[42][0],vnu_pa_msg[41][0],vnu_pa_msg[40][0],vnu_pa_msg[39][0],vnu_pa_msg[38][0],vnu_pa_msg[37][0],vnu_pa_msg[36][0],vnu_pa_msg[35][0],vnu_pa_msg[34][0],vnu_pa_msg[33][0],vnu_pa_msg[32][0],vnu_pa_msg[31][0],vnu_pa_msg[30][0],vnu_pa_msg[29][0],vnu_pa_msg[28][0],vnu_pa_msg[27][0],vnu_pa_msg[26][0],vnu_pa_msg[25][0],vnu_pa_msg[24][0],vnu_pa_msg[23][0],vnu_pa_msg[22][0],vnu_pa_msg[21][0],vnu_pa_msg[20][0],vnu_pa_msg[19][0],vnu_pa_msg[18][0],vnu_pa_msg[17][0],vnu_pa_msg[16][0],vnu_pa_msg[15][0],vnu_pa_msg[14][0],vnu_pa_msg[13][0],vnu_pa_msg[12][0],vnu_pa_msg[11][0],vnu_pa_msg[10][0],vnu_pa_msg[9][0],vnu_pa_msg[8][0],vnu_pa_msg[7][0],vnu_pa_msg[6][0],vnu_pa_msg[5][0],vnu_pa_msg[4][0],vnu_pa_msg[3][0],vnu_pa_msg[2][0],vnu_pa_msg[1][0],vnu_pa_msg[0][0]};
assign pa_to_ch_ram[CH_DATA_WIDTH-1:0] = {vnu_pa_msg[84][QUAN_SIZE-1:0],vnu_pa_msg[83][QUAN_SIZE-1:0],vnu_pa_msg[82][QUAN_SIZE-1:0],vnu_pa_msg[81][QUAN_SIZE-1:0],vnu_pa_msg[80][QUAN_SIZE-1:0],vnu_pa_msg[79][QUAN_SIZE-1:0],vnu_pa_msg[78][QUAN_SIZE-1:0],vnu_pa_msg[77][QUAN_SIZE-1:0],vnu_pa_msg[76][QUAN_SIZE-1:0],vnu_pa_msg[75][QUAN_SIZE-1:0],vnu_pa_msg[74][QUAN_SIZE-1:0],vnu_pa_msg[73][QUAN_SIZE-1:0],vnu_pa_msg[72][QUAN_SIZE-1:0],vnu_pa_msg[71][QUAN_SIZE-1:0],vnu_pa_msg[70][QUAN_SIZE-1:0],vnu_pa_msg[69][QUAN_SIZE-1:0],vnu_pa_msg[68][QUAN_SIZE-1:0],vnu_pa_msg[67][QUAN_SIZE-1:0],vnu_pa_msg[66][QUAN_SIZE-1:0],vnu_pa_msg[65][QUAN_SIZE-1:0],vnu_pa_msg[64][QUAN_SIZE-1:0],vnu_pa_msg[63][QUAN_SIZE-1:0],vnu_pa_msg[62][QUAN_SIZE-1:0],vnu_pa_msg[61][QUAN_SIZE-1:0],vnu_pa_msg[60][QUAN_SIZE-1:0],vnu_pa_msg[59][QUAN_SIZE-1:0],vnu_pa_msg[58][QUAN_SIZE-1:0],vnu_pa_msg[57][QUAN_SIZE-1:0],vnu_pa_msg[56][QUAN_SIZE-1:0],vnu_pa_msg[55][QUAN_SIZE-1:0],vnu_pa_msg[54][QUAN_SIZE-1:0],vnu_pa_msg[53][QUAN_SIZE-1:0],vnu_pa_msg[52][QUAN_SIZE-1:0],vnu_pa_msg[51][QUAN_SIZE-1:0],vnu_pa_msg[50][QUAN_SIZE-1:0],vnu_pa_msg[49][QUAN_SIZE-1:0],vnu_pa_msg[48][QUAN_SIZE-1:0],vnu_pa_msg[47][QUAN_SIZE-1:0],vnu_pa_msg[46][QUAN_SIZE-1:0],vnu_pa_msg[45][QUAN_SIZE-1:0],vnu_pa_msg[44][QUAN_SIZE-1:0],vnu_pa_msg[43][QUAN_SIZE-1:0],vnu_pa_msg[42][QUAN_SIZE-1:0],vnu_pa_msg[41][QUAN_SIZE-1:0],vnu_pa_msg[40][QUAN_SIZE-1:0],vnu_pa_msg[39][QUAN_SIZE-1:0],vnu_pa_msg[38][QUAN_SIZE-1:0],vnu_pa_msg[37][QUAN_SIZE-1:0],vnu_pa_msg[36][QUAN_SIZE-1:0],vnu_pa_msg[35][QUAN_SIZE-1:0],vnu_pa_msg[34][QUAN_SIZE-1:0],vnu_pa_msg[33][QUAN_SIZE-1:0],vnu_pa_msg[32][QUAN_SIZE-1:0],vnu_pa_msg[31][QUAN_SIZE-1:0],vnu_pa_msg[30][QUAN_SIZE-1:0],vnu_pa_msg[29][QUAN_SIZE-1:0],vnu_pa_msg[28][QUAN_SIZE-1:0],vnu_pa_msg[27][QUAN_SIZE-1:0],vnu_pa_msg[26][QUAN_SIZE-1:0],vnu_pa_msg[25][QUAN_SIZE-1:0],vnu_pa_msg[24][QUAN_SIZE-1:0],vnu_pa_msg[23][QUAN_SIZE-1:0],vnu_pa_msg[22][QUAN_SIZE-1:0],vnu_pa_msg[21][QUAN_SIZE-1:0],vnu_pa_msg[20][QUAN_SIZE-1:0],vnu_pa_msg[19][QUAN_SIZE-1:0],vnu_pa_msg[18][QUAN_SIZE-1:0],vnu_pa_msg[17][QUAN_SIZE-1:0],vnu_pa_msg[16][QUAN_SIZE-1:0],vnu_pa_msg[15][QUAN_SIZE-1:0],vnu_pa_msg[14][QUAN_SIZE-1:0],vnu_pa_msg[13][QUAN_SIZE-1:0],vnu_pa_msg[12][QUAN_SIZE-1:0],vnu_pa_msg[11][QUAN_SIZE-1:0],vnu_pa_msg[10][QUAN_SIZE-1:0],vnu_pa_msg[9][QUAN_SIZE-1:0],vnu_pa_msg[8][QUAN_SIZE-1:0],vnu_pa_msg[7][QUAN_SIZE-1:0],vnu_pa_msg[6][QUAN_SIZE-1:0],vnu_pa_msg[5][QUAN_SIZE-1:0],vnu_pa_msg[4][QUAN_SIZE-1:0],vnu_pa_msg[3][QUAN_SIZE-1:0],vnu_pa_msg[2][QUAN_SIZE-1:0],vnu_pa_msg[1][QUAN_SIZE-1:0],vnu_pa_msg[0][QUAN_SIZE-1:0]};
endmodule
`endif