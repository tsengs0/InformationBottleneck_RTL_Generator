`include "define.vh"

module top_layer_decoder (

);


endmodule