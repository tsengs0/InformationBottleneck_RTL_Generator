module ib_proc_wrapper #(
	parameter CN_ROM_RD_BW = 6,
	parameter CN_ROM_ADDR_BW = 10,
	parameter CN_PAGE_ADDR_BW = 5,
	parameter CN_DEGREE = 6,
	parameter IB_CNU_DECOMP_funNum = 4,
	parameter CN_NUM = 102,
	parameter CNU6_INSTANTIATE_NUM = 51,
	parameter CNU6_INSTANTIATE_UNIT = 2,

	parameter VN_ROM_RD_BW = 8,
	parameter VN_ROM_ADDR_BW = 11,
	parameter VN_PAGE_ADDR_BW = 6,
	parameter DN_ROM_RD_BW = 8,
	parameter DN_ROM_ADDR_BW = 11,
	parameter DN_PAGE_ADDR_BW = 6,
	parameter VN_DEGREE = 3,
	parameter IB_VNU_DECOMP_funNum = 2,
	parameter VN_NUM = 204,
	parameter VNU3_INSTANTIATE_NUM = 51,
	parameter VNU3_INSTANTIATE_UNIT = 4,
	parameter QUAN_SIZE = 4,
	parameter MSG_WIDTH = 4,
	parameter DATAPATH_WIDTH = 4
) (
	output wire [VN_NUM-1:0] hard_decision,

	input wire [DATAPATH_WIDTH-1:0] ch_msg_0,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_1,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_2,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_3,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_4,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_5,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_6,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_7,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_8,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_9,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_10,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_11,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_12,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_13,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_14,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_15,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_16,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_17,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_18,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_19,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_20,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_21,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_22,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_23,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_24,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_25,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_26,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_27,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_28,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_29,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_30,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_31,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_32,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_33,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_34,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_35,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_36,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_37,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_38,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_39,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_40,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_41,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_42,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_43,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_44,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_45,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_46,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_47,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_48,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_49,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_50,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_51,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_52,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_53,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_54,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_55,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_56,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_57,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_58,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_59,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_60,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_61,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_62,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_63,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_64,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_65,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_66,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_67,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_68,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_69,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_70,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_71,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_72,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_73,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_74,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_75,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_76,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_77,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_78,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_79,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_80,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_81,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_82,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_83,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_84,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_85,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_86,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_87,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_88,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_89,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_90,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_91,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_92,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_93,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_94,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_95,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_96,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_97,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_98,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_99,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_100,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_101,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_102,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_103,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_104,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_105,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_106,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_107,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_108,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_109,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_110,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_111,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_112,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_113,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_114,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_115,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_116,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_117,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_118,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_119,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_120,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_121,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_122,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_123,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_124,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_125,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_126,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_127,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_128,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_129,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_130,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_131,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_132,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_133,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_134,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_135,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_136,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_137,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_138,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_139,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_140,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_141,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_142,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_143,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_144,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_145,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_146,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_147,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_148,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_149,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_150,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_151,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_152,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_153,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_154,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_155,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_156,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_157,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_158,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_159,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_160,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_161,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_162,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_163,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_164,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_165,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_166,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_167,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_168,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_169,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_170,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_171,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_172,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_173,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_174,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_175,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_176,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_177,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_178,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_179,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_180,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_181,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_182,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_183,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_184,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_185,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_186,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_187,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_188,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_189,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_190,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_191,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_192,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_193,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_194,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_195,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_196,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_197,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_198,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_199,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_200,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_201,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_202,
	input wire [DATAPATH_WIDTH-1:0] ch_msg_203,
	input wire read_clk,
	input wire cnu_read_addr_offset,
	input wire vnu_read_addr_offset,
	input wire v2c_latch_en,
	input wire c2v_latch_en,
	input wire v2c_src,
	input wire [1:0] parallel_en,
	input wire [1:0] load,

	// Iteration-Refresh Page Address
	input wire [CN_PAGE_ADDR_BW+1-1:0] cnu_page_addr_ram_0, // the MSB decides refreshed target, i.e., upper page group or lower page group
	input wire [CN_PAGE_ADDR_BW+1-1:0] cnu_page_addr_ram_1, // the MSB decides refreshed target, i.e., upper page group or lower page group
	input wire [CN_PAGE_ADDR_BW+1-1:0] cnu_page_addr_ram_2, // the MSB decides refreshed target, i.e., upper page group or lower page group
	input wire [CN_PAGE_ADDR_BW+1-1:0] cnu_page_addr_ram_3, // the MSB decides refreshed target, i.e., upper page group or lower page group
	input wire [VN_PAGE_ADDR_BW+1-1:0] vnu_page_addr_ram_0, // the MSB decides refreshed target, i.e., upper page group or lower page group
	input wire [VN_PAGE_ADDR_BW+1-1:0] vnu_page_addr_ram_1, // the MSB decides refreshed target, i.e., upper page group or lower page group
	input wire [VN_PAGE_ADDR_BW+1-1:0] vnu_page_addr_ram_2, // the MSB decides refreshed target, i.e., upper page group or lower page group // the last one is for decision node
	//Iteration-Refresh Page Data
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataA_0, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataB_0, // from portB of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataA_1, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataB_1, // from portB of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataA_2, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataB_2, // from portB of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataA_3, // from portA of IB-ROM
	input wire [CN_ROM_RD_BW-1:0] cnu_ram_write_dataB_3, // from portB of IB-ROM
	input wire [VN_ROM_RD_BW-1:0] vnu_ram_write_dataA_0, // from portA of IB-ROM
	input wire [VN_ROM_RD_BW-1:0] vnu_ram_write_dataB_0, // from portB of IB-ROM
	input wire [VN_ROM_RD_BW-1:0] vnu_ram_write_dataA_1, // from portA of IB-ROM
	input wire [VN_ROM_RD_BW-1:0] vnu_ram_write_dataB_1, // from portB of IB-ROM
	input wire [DN_ROM_RD_BW-1:0] vnu_ram_write_dataA_2, // from portA of IB-ROM (for decision node)
	input wire [DN_ROM_RD_BW-1:0] vnu_ram_write_dataB_2, // from portB of IB-ROM (for decision node)

	input wire [3:0] cnu_ib_ram_we,
	input wire [2:0] vnu_ib_ram_we,
	input wire cn_write_clk,
	input wire vn_write_clk,
	input wire dn_write_clk
);

// Net-type interfaces (direction is RouteNetworkModule-centric)
//        -------
//       |  cnu  |
//        -------
//         |  ^        
// c2v_in  |  | v2c_out
//         v  |        
//       ----------
//      |   Route  |
//      | __    __ |
//      |   \  /   |
//      |    \/    |
//      |    /\    |
//      | __/  \__ |
//       -----------
//          |  ^       
// c2v_out  |  | v2c_in
//          v  |       
//         -------
//        |  vnu  |
//         -------
wire [DATAPATH_WIDTH-1:0] c2v_in0 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] v2c_out0 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_in1 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] v2c_out1 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_in2 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] v2c_out2 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_in3 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] v2c_out3 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_in4 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] v2c_out4 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_in5 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] v2c_out5 [0:CN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_out0 [0:VN_NUM-1]; 
wire [DATAPATH_WIDTH-1:0] v2c_in0 [0:VN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_out1 [0:VN_NUM-1]; 
wire [DATAPATH_WIDTH-1:0] v2c_in1 [0:VN_NUM-1];
wire [DATAPATH_WIDTH-1:0] c2v_out2 [0:VN_NUM-1]; 
wire [DATAPATH_WIDTH-1:0] v2c_in2 [0:VN_NUM-1];

// Instantiation of CNU IB-RAM wrapper
cnu6_ib_ram_wrapper #(
	.CN_ROM_RD_BW          (CN_ROM_RD_BW         ),
	.CN_ROM_ADDR_BW        (CN_ROM_ADDR_BW       ),
	.CN_PAGE_ADDR_BW       (CN_PAGE_ADDR_BW      ),
	.CN_DEGREE	          (CN_DEGREE            ),
	.IB_CNU_DECOMP_funNum  (IB_CNU_DECOMP_funNum ),
	.CN_NUM                (CN_NUM               ),
	.CNU6_INSTANTIATE_NUM  (CNU6_INSTANTIATE_NUM ),
	.CNU6_INSTANTIATE_UNIT (CNU6_INSTANTIATE_UNIT),
	.QUAN_SIZE             (QUAN_SIZE            ),
	.DATAPATH_WIDTH        (DATAPATH_WIDTH       )
) cnu_ib_ram_wrapper_u0 (
	.c2v_0_out0(c2v_in0[0]),
	.c2v_0_out1(c2v_in1[0]),
	.c2v_0_out2(c2v_in2[0]),
	.c2v_0_out3(c2v_in3[0]),
	.c2v_0_out4(c2v_in4[0]),
	.c2v_0_out5(c2v_in5[0]),
	.c2v_1_out0(c2v_in0[1]),
	.c2v_1_out1(c2v_in1[1]),
	.c2v_1_out2(c2v_in2[1]),
	.c2v_1_out3(c2v_in3[1]),
	.c2v_1_out4(c2v_in4[1]),
	.c2v_1_out5(c2v_in5[1]),
	.c2v_2_out0(c2v_in0[2]),
	.c2v_2_out1(c2v_in1[2]),
	.c2v_2_out2(c2v_in2[2]),
	.c2v_2_out3(c2v_in3[2]),
	.c2v_2_out4(c2v_in4[2]),
	.c2v_2_out5(c2v_in5[2]),
	.c2v_3_out0(c2v_in0[3]),
	.c2v_3_out1(c2v_in1[3]),
	.c2v_3_out2(c2v_in2[3]),
	.c2v_3_out3(c2v_in3[3]),
	.c2v_3_out4(c2v_in4[3]),
	.c2v_3_out5(c2v_in5[3]),
	.c2v_4_out0(c2v_in0[4]),
	.c2v_4_out1(c2v_in1[4]),
	.c2v_4_out2(c2v_in2[4]),
	.c2v_4_out3(c2v_in3[4]),
	.c2v_4_out4(c2v_in4[4]),
	.c2v_4_out5(c2v_in5[4]),
	.c2v_5_out0(c2v_in0[5]),
	.c2v_5_out1(c2v_in1[5]),
	.c2v_5_out2(c2v_in2[5]),
	.c2v_5_out3(c2v_in3[5]),
	.c2v_5_out4(c2v_in4[5]),
	.c2v_5_out5(c2v_in5[5]),
	.c2v_6_out0(c2v_in0[6]),
	.c2v_6_out1(c2v_in1[6]),
	.c2v_6_out2(c2v_in2[6]),
	.c2v_6_out3(c2v_in3[6]),
	.c2v_6_out4(c2v_in4[6]),
	.c2v_6_out5(c2v_in5[6]),
	.c2v_7_out0(c2v_in0[7]),
	.c2v_7_out1(c2v_in1[7]),
	.c2v_7_out2(c2v_in2[7]),
	.c2v_7_out3(c2v_in3[7]),
	.c2v_7_out4(c2v_in4[7]),
	.c2v_7_out5(c2v_in5[7]),
	.c2v_8_out0(c2v_in0[8]),
	.c2v_8_out1(c2v_in1[8]),
	.c2v_8_out2(c2v_in2[8]),
	.c2v_8_out3(c2v_in3[8]),
	.c2v_8_out4(c2v_in4[8]),
	.c2v_8_out5(c2v_in5[8]),
	.c2v_9_out0(c2v_in0[9]),
	.c2v_9_out1(c2v_in1[9]),
	.c2v_9_out2(c2v_in2[9]),
	.c2v_9_out3(c2v_in3[9]),
	.c2v_9_out4(c2v_in4[9]),
	.c2v_9_out5(c2v_in5[9]),
	.c2v_10_out0(c2v_in0[10]),
	.c2v_10_out1(c2v_in1[10]),
	.c2v_10_out2(c2v_in2[10]),
	.c2v_10_out3(c2v_in3[10]),
	.c2v_10_out4(c2v_in4[10]),
	.c2v_10_out5(c2v_in5[10]),
	.c2v_11_out0(c2v_in0[11]),
	.c2v_11_out1(c2v_in1[11]),
	.c2v_11_out2(c2v_in2[11]),
	.c2v_11_out3(c2v_in3[11]),
	.c2v_11_out4(c2v_in4[11]),
	.c2v_11_out5(c2v_in5[11]),
	.c2v_12_out0(c2v_in0[12]),
	.c2v_12_out1(c2v_in1[12]),
	.c2v_12_out2(c2v_in2[12]),
	.c2v_12_out3(c2v_in3[12]),
	.c2v_12_out4(c2v_in4[12]),
	.c2v_12_out5(c2v_in5[12]),
	.c2v_13_out0(c2v_in0[13]),
	.c2v_13_out1(c2v_in1[13]),
	.c2v_13_out2(c2v_in2[13]),
	.c2v_13_out3(c2v_in3[13]),
	.c2v_13_out4(c2v_in4[13]),
	.c2v_13_out5(c2v_in5[13]),
	.c2v_14_out0(c2v_in0[14]),
	.c2v_14_out1(c2v_in1[14]),
	.c2v_14_out2(c2v_in2[14]),
	.c2v_14_out3(c2v_in3[14]),
	.c2v_14_out4(c2v_in4[14]),
	.c2v_14_out5(c2v_in5[14]),
	.c2v_15_out0(c2v_in0[15]),
	.c2v_15_out1(c2v_in1[15]),
	.c2v_15_out2(c2v_in2[15]),
	.c2v_15_out3(c2v_in3[15]),
	.c2v_15_out4(c2v_in4[15]),
	.c2v_15_out5(c2v_in5[15]),
	.c2v_16_out0(c2v_in0[16]),
	.c2v_16_out1(c2v_in1[16]),
	.c2v_16_out2(c2v_in2[16]),
	.c2v_16_out3(c2v_in3[16]),
	.c2v_16_out4(c2v_in4[16]),
	.c2v_16_out5(c2v_in5[16]),
	.c2v_17_out0(c2v_in0[17]),
	.c2v_17_out1(c2v_in1[17]),
	.c2v_17_out2(c2v_in2[17]),
	.c2v_17_out3(c2v_in3[17]),
	.c2v_17_out4(c2v_in4[17]),
	.c2v_17_out5(c2v_in5[17]),
	.c2v_18_out0(c2v_in0[18]),
	.c2v_18_out1(c2v_in1[18]),
	.c2v_18_out2(c2v_in2[18]),
	.c2v_18_out3(c2v_in3[18]),
	.c2v_18_out4(c2v_in4[18]),
	.c2v_18_out5(c2v_in5[18]),
	.c2v_19_out0(c2v_in0[19]),
	.c2v_19_out1(c2v_in1[19]),
	.c2v_19_out2(c2v_in2[19]),
	.c2v_19_out3(c2v_in3[19]),
	.c2v_19_out4(c2v_in4[19]),
	.c2v_19_out5(c2v_in5[19]),
	.c2v_20_out0(c2v_in0[20]),
	.c2v_20_out1(c2v_in1[20]),
	.c2v_20_out2(c2v_in2[20]),
	.c2v_20_out3(c2v_in3[20]),
	.c2v_20_out4(c2v_in4[20]),
	.c2v_20_out5(c2v_in5[20]),
	.c2v_21_out0(c2v_in0[21]),
	.c2v_21_out1(c2v_in1[21]),
	.c2v_21_out2(c2v_in2[21]),
	.c2v_21_out3(c2v_in3[21]),
	.c2v_21_out4(c2v_in4[21]),
	.c2v_21_out5(c2v_in5[21]),
	.c2v_22_out0(c2v_in0[22]),
	.c2v_22_out1(c2v_in1[22]),
	.c2v_22_out2(c2v_in2[22]),
	.c2v_22_out3(c2v_in3[22]),
	.c2v_22_out4(c2v_in4[22]),
	.c2v_22_out5(c2v_in5[22]),
	.c2v_23_out0(c2v_in0[23]),
	.c2v_23_out1(c2v_in1[23]),
	.c2v_23_out2(c2v_in2[23]),
	.c2v_23_out3(c2v_in3[23]),
	.c2v_23_out4(c2v_in4[23]),
	.c2v_23_out5(c2v_in5[23]),
	.c2v_24_out0(c2v_in0[24]),
	.c2v_24_out1(c2v_in1[24]),
	.c2v_24_out2(c2v_in2[24]),
	.c2v_24_out3(c2v_in3[24]),
	.c2v_24_out4(c2v_in4[24]),
	.c2v_24_out5(c2v_in5[24]),
	.c2v_25_out0(c2v_in0[25]),
	.c2v_25_out1(c2v_in1[25]),
	.c2v_25_out2(c2v_in2[25]),
	.c2v_25_out3(c2v_in3[25]),
	.c2v_25_out4(c2v_in4[25]),
	.c2v_25_out5(c2v_in5[25]),
	.c2v_26_out0(c2v_in0[26]),
	.c2v_26_out1(c2v_in1[26]),
	.c2v_26_out2(c2v_in2[26]),
	.c2v_26_out3(c2v_in3[26]),
	.c2v_26_out4(c2v_in4[26]),
	.c2v_26_out5(c2v_in5[26]),
	.c2v_27_out0(c2v_in0[27]),
	.c2v_27_out1(c2v_in1[27]),
	.c2v_27_out2(c2v_in2[27]),
	.c2v_27_out3(c2v_in3[27]),
	.c2v_27_out4(c2v_in4[27]),
	.c2v_27_out5(c2v_in5[27]),
	.c2v_28_out0(c2v_in0[28]),
	.c2v_28_out1(c2v_in1[28]),
	.c2v_28_out2(c2v_in2[28]),
	.c2v_28_out3(c2v_in3[28]),
	.c2v_28_out4(c2v_in4[28]),
	.c2v_28_out5(c2v_in5[28]),
	.c2v_29_out0(c2v_in0[29]),
	.c2v_29_out1(c2v_in1[29]),
	.c2v_29_out2(c2v_in2[29]),
	.c2v_29_out3(c2v_in3[29]),
	.c2v_29_out4(c2v_in4[29]),
	.c2v_29_out5(c2v_in5[29]),
	.c2v_30_out0(c2v_in0[30]),
	.c2v_30_out1(c2v_in1[30]),
	.c2v_30_out2(c2v_in2[30]),
	.c2v_30_out3(c2v_in3[30]),
	.c2v_30_out4(c2v_in4[30]),
	.c2v_30_out5(c2v_in5[30]),
	.c2v_31_out0(c2v_in0[31]),
	.c2v_31_out1(c2v_in1[31]),
	.c2v_31_out2(c2v_in2[31]),
	.c2v_31_out3(c2v_in3[31]),
	.c2v_31_out4(c2v_in4[31]),
	.c2v_31_out5(c2v_in5[31]),
	.c2v_32_out0(c2v_in0[32]),
	.c2v_32_out1(c2v_in1[32]),
	.c2v_32_out2(c2v_in2[32]),
	.c2v_32_out3(c2v_in3[32]),
	.c2v_32_out4(c2v_in4[32]),
	.c2v_32_out5(c2v_in5[32]),
	.c2v_33_out0(c2v_in0[33]),
	.c2v_33_out1(c2v_in1[33]),
	.c2v_33_out2(c2v_in2[33]),
	.c2v_33_out3(c2v_in3[33]),
	.c2v_33_out4(c2v_in4[33]),
	.c2v_33_out5(c2v_in5[33]),
	.c2v_34_out0(c2v_in0[34]),
	.c2v_34_out1(c2v_in1[34]),
	.c2v_34_out2(c2v_in2[34]),
	.c2v_34_out3(c2v_in3[34]),
	.c2v_34_out4(c2v_in4[34]),
	.c2v_34_out5(c2v_in5[34]),
	.c2v_35_out0(c2v_in0[35]),
	.c2v_35_out1(c2v_in1[35]),
	.c2v_35_out2(c2v_in2[35]),
	.c2v_35_out3(c2v_in3[35]),
	.c2v_35_out4(c2v_in4[35]),
	.c2v_35_out5(c2v_in5[35]),
	.c2v_36_out0(c2v_in0[36]),
	.c2v_36_out1(c2v_in1[36]),
	.c2v_36_out2(c2v_in2[36]),
	.c2v_36_out3(c2v_in3[36]),
	.c2v_36_out4(c2v_in4[36]),
	.c2v_36_out5(c2v_in5[36]),
	.c2v_37_out0(c2v_in0[37]),
	.c2v_37_out1(c2v_in1[37]),
	.c2v_37_out2(c2v_in2[37]),
	.c2v_37_out3(c2v_in3[37]),
	.c2v_37_out4(c2v_in4[37]),
	.c2v_37_out5(c2v_in5[37]),
	.c2v_38_out0(c2v_in0[38]),
	.c2v_38_out1(c2v_in1[38]),
	.c2v_38_out2(c2v_in2[38]),
	.c2v_38_out3(c2v_in3[38]),
	.c2v_38_out4(c2v_in4[38]),
	.c2v_38_out5(c2v_in5[38]),
	.c2v_39_out0(c2v_in0[39]),
	.c2v_39_out1(c2v_in1[39]),
	.c2v_39_out2(c2v_in2[39]),
	.c2v_39_out3(c2v_in3[39]),
	.c2v_39_out4(c2v_in4[39]),
	.c2v_39_out5(c2v_in5[39]),
	.c2v_40_out0(c2v_in0[40]),
	.c2v_40_out1(c2v_in1[40]),
	.c2v_40_out2(c2v_in2[40]),
	.c2v_40_out3(c2v_in3[40]),
	.c2v_40_out4(c2v_in4[40]),
	.c2v_40_out5(c2v_in5[40]),
	.c2v_41_out0(c2v_in0[41]),
	.c2v_41_out1(c2v_in1[41]),
	.c2v_41_out2(c2v_in2[41]),
	.c2v_41_out3(c2v_in3[41]),
	.c2v_41_out4(c2v_in4[41]),
	.c2v_41_out5(c2v_in5[41]),
	.c2v_42_out0(c2v_in0[42]),
	.c2v_42_out1(c2v_in1[42]),
	.c2v_42_out2(c2v_in2[42]),
	.c2v_42_out3(c2v_in3[42]),
	.c2v_42_out4(c2v_in4[42]),
	.c2v_42_out5(c2v_in5[42]),
	.c2v_43_out0(c2v_in0[43]),
	.c2v_43_out1(c2v_in1[43]),
	.c2v_43_out2(c2v_in2[43]),
	.c2v_43_out3(c2v_in3[43]),
	.c2v_43_out4(c2v_in4[43]),
	.c2v_43_out5(c2v_in5[43]),
	.c2v_44_out0(c2v_in0[44]),
	.c2v_44_out1(c2v_in1[44]),
	.c2v_44_out2(c2v_in2[44]),
	.c2v_44_out3(c2v_in3[44]),
	.c2v_44_out4(c2v_in4[44]),
	.c2v_44_out5(c2v_in5[44]),
	.c2v_45_out0(c2v_in0[45]),
	.c2v_45_out1(c2v_in1[45]),
	.c2v_45_out2(c2v_in2[45]),
	.c2v_45_out3(c2v_in3[45]),
	.c2v_45_out4(c2v_in4[45]),
	.c2v_45_out5(c2v_in5[45]),
	.c2v_46_out0(c2v_in0[46]),
	.c2v_46_out1(c2v_in1[46]),
	.c2v_46_out2(c2v_in2[46]),
	.c2v_46_out3(c2v_in3[46]),
	.c2v_46_out4(c2v_in4[46]),
	.c2v_46_out5(c2v_in5[46]),
	.c2v_47_out0(c2v_in0[47]),
	.c2v_47_out1(c2v_in1[47]),
	.c2v_47_out2(c2v_in2[47]),
	.c2v_47_out3(c2v_in3[47]),
	.c2v_47_out4(c2v_in4[47]),
	.c2v_47_out5(c2v_in5[47]),
	.c2v_48_out0(c2v_in0[48]),
	.c2v_48_out1(c2v_in1[48]),
	.c2v_48_out2(c2v_in2[48]),
	.c2v_48_out3(c2v_in3[48]),
	.c2v_48_out4(c2v_in4[48]),
	.c2v_48_out5(c2v_in5[48]),
	.c2v_49_out0(c2v_in0[49]),
	.c2v_49_out1(c2v_in1[49]),
	.c2v_49_out2(c2v_in2[49]),
	.c2v_49_out3(c2v_in3[49]),
	.c2v_49_out4(c2v_in4[49]),
	.c2v_49_out5(c2v_in5[49]),
	.c2v_50_out0(c2v_in0[50]),
	.c2v_50_out1(c2v_in1[50]),
	.c2v_50_out2(c2v_in2[50]),
	.c2v_50_out3(c2v_in3[50]),
	.c2v_50_out4(c2v_in4[50]),
	.c2v_50_out5(c2v_in5[50]),
	.c2v_51_out0(c2v_in0[51]),
	.c2v_51_out1(c2v_in1[51]),
	.c2v_51_out2(c2v_in2[51]),
	.c2v_51_out3(c2v_in3[51]),
	.c2v_51_out4(c2v_in4[51]),
	.c2v_51_out5(c2v_in5[51]),
	.c2v_52_out0(c2v_in0[52]),
	.c2v_52_out1(c2v_in1[52]),
	.c2v_52_out2(c2v_in2[52]),
	.c2v_52_out3(c2v_in3[52]),
	.c2v_52_out4(c2v_in4[52]),
	.c2v_52_out5(c2v_in5[52]),
	.c2v_53_out0(c2v_in0[53]),
	.c2v_53_out1(c2v_in1[53]),
	.c2v_53_out2(c2v_in2[53]),
	.c2v_53_out3(c2v_in3[53]),
	.c2v_53_out4(c2v_in4[53]),
	.c2v_53_out5(c2v_in5[53]),
	.c2v_54_out0(c2v_in0[54]),
	.c2v_54_out1(c2v_in1[54]),
	.c2v_54_out2(c2v_in2[54]),
	.c2v_54_out3(c2v_in3[54]),
	.c2v_54_out4(c2v_in4[54]),
	.c2v_54_out5(c2v_in5[54]),
	.c2v_55_out0(c2v_in0[55]),
	.c2v_55_out1(c2v_in1[55]),
	.c2v_55_out2(c2v_in2[55]),
	.c2v_55_out3(c2v_in3[55]),
	.c2v_55_out4(c2v_in4[55]),
	.c2v_55_out5(c2v_in5[55]),
	.c2v_56_out0(c2v_in0[56]),
	.c2v_56_out1(c2v_in1[56]),
	.c2v_56_out2(c2v_in2[56]),
	.c2v_56_out3(c2v_in3[56]),
	.c2v_56_out4(c2v_in4[56]),
	.c2v_56_out5(c2v_in5[56]),
	.c2v_57_out0(c2v_in0[57]),
	.c2v_57_out1(c2v_in1[57]),
	.c2v_57_out2(c2v_in2[57]),
	.c2v_57_out3(c2v_in3[57]),
	.c2v_57_out4(c2v_in4[57]),
	.c2v_57_out5(c2v_in5[57]),
	.c2v_58_out0(c2v_in0[58]),
	.c2v_58_out1(c2v_in1[58]),
	.c2v_58_out2(c2v_in2[58]),
	.c2v_58_out3(c2v_in3[58]),
	.c2v_58_out4(c2v_in4[58]),
	.c2v_58_out5(c2v_in5[58]),
	.c2v_59_out0(c2v_in0[59]),
	.c2v_59_out1(c2v_in1[59]),
	.c2v_59_out2(c2v_in2[59]),
	.c2v_59_out3(c2v_in3[59]),
	.c2v_59_out4(c2v_in4[59]),
	.c2v_59_out5(c2v_in5[59]),
	.c2v_60_out0(c2v_in0[60]),
	.c2v_60_out1(c2v_in1[60]),
	.c2v_60_out2(c2v_in2[60]),
	.c2v_60_out3(c2v_in3[60]),
	.c2v_60_out4(c2v_in4[60]),
	.c2v_60_out5(c2v_in5[60]),
	.c2v_61_out0(c2v_in0[61]),
	.c2v_61_out1(c2v_in1[61]),
	.c2v_61_out2(c2v_in2[61]),
	.c2v_61_out3(c2v_in3[61]),
	.c2v_61_out4(c2v_in4[61]),
	.c2v_61_out5(c2v_in5[61]),
	.c2v_62_out0(c2v_in0[62]),
	.c2v_62_out1(c2v_in1[62]),
	.c2v_62_out2(c2v_in2[62]),
	.c2v_62_out3(c2v_in3[62]),
	.c2v_62_out4(c2v_in4[62]),
	.c2v_62_out5(c2v_in5[62]),
	.c2v_63_out0(c2v_in0[63]),
	.c2v_63_out1(c2v_in1[63]),
	.c2v_63_out2(c2v_in2[63]),
	.c2v_63_out3(c2v_in3[63]),
	.c2v_63_out4(c2v_in4[63]),
	.c2v_63_out5(c2v_in5[63]),
	.c2v_64_out0(c2v_in0[64]),
	.c2v_64_out1(c2v_in1[64]),
	.c2v_64_out2(c2v_in2[64]),
	.c2v_64_out3(c2v_in3[64]),
	.c2v_64_out4(c2v_in4[64]),
	.c2v_64_out5(c2v_in5[64]),
	.c2v_65_out0(c2v_in0[65]),
	.c2v_65_out1(c2v_in1[65]),
	.c2v_65_out2(c2v_in2[65]),
	.c2v_65_out3(c2v_in3[65]),
	.c2v_65_out4(c2v_in4[65]),
	.c2v_65_out5(c2v_in5[65]),
	.c2v_66_out0(c2v_in0[66]),
	.c2v_66_out1(c2v_in1[66]),
	.c2v_66_out2(c2v_in2[66]),
	.c2v_66_out3(c2v_in3[66]),
	.c2v_66_out4(c2v_in4[66]),
	.c2v_66_out5(c2v_in5[66]),
	.c2v_67_out0(c2v_in0[67]),
	.c2v_67_out1(c2v_in1[67]),
	.c2v_67_out2(c2v_in2[67]),
	.c2v_67_out3(c2v_in3[67]),
	.c2v_67_out4(c2v_in4[67]),
	.c2v_67_out5(c2v_in5[67]),
	.c2v_68_out0(c2v_in0[68]),
	.c2v_68_out1(c2v_in1[68]),
	.c2v_68_out2(c2v_in2[68]),
	.c2v_68_out3(c2v_in3[68]),
	.c2v_68_out4(c2v_in4[68]),
	.c2v_68_out5(c2v_in5[68]),
	.c2v_69_out0(c2v_in0[69]),
	.c2v_69_out1(c2v_in1[69]),
	.c2v_69_out2(c2v_in2[69]),
	.c2v_69_out3(c2v_in3[69]),
	.c2v_69_out4(c2v_in4[69]),
	.c2v_69_out5(c2v_in5[69]),
	.c2v_70_out0(c2v_in0[70]),
	.c2v_70_out1(c2v_in1[70]),
	.c2v_70_out2(c2v_in2[70]),
	.c2v_70_out3(c2v_in3[70]),
	.c2v_70_out4(c2v_in4[70]),
	.c2v_70_out5(c2v_in5[70]),
	.c2v_71_out0(c2v_in0[71]),
	.c2v_71_out1(c2v_in1[71]),
	.c2v_71_out2(c2v_in2[71]),
	.c2v_71_out3(c2v_in3[71]),
	.c2v_71_out4(c2v_in4[71]),
	.c2v_71_out5(c2v_in5[71]),
	.c2v_72_out0(c2v_in0[72]),
	.c2v_72_out1(c2v_in1[72]),
	.c2v_72_out2(c2v_in2[72]),
	.c2v_72_out3(c2v_in3[72]),
	.c2v_72_out4(c2v_in4[72]),
	.c2v_72_out5(c2v_in5[72]),
	.c2v_73_out0(c2v_in0[73]),
	.c2v_73_out1(c2v_in1[73]),
	.c2v_73_out2(c2v_in2[73]),
	.c2v_73_out3(c2v_in3[73]),
	.c2v_73_out4(c2v_in4[73]),
	.c2v_73_out5(c2v_in5[73]),
	.c2v_74_out0(c2v_in0[74]),
	.c2v_74_out1(c2v_in1[74]),
	.c2v_74_out2(c2v_in2[74]),
	.c2v_74_out3(c2v_in3[74]),
	.c2v_74_out4(c2v_in4[74]),
	.c2v_74_out5(c2v_in5[74]),
	.c2v_75_out0(c2v_in0[75]),
	.c2v_75_out1(c2v_in1[75]),
	.c2v_75_out2(c2v_in2[75]),
	.c2v_75_out3(c2v_in3[75]),
	.c2v_75_out4(c2v_in4[75]),
	.c2v_75_out5(c2v_in5[75]),
	.c2v_76_out0(c2v_in0[76]),
	.c2v_76_out1(c2v_in1[76]),
	.c2v_76_out2(c2v_in2[76]),
	.c2v_76_out3(c2v_in3[76]),
	.c2v_76_out4(c2v_in4[76]),
	.c2v_76_out5(c2v_in5[76]),
	.c2v_77_out0(c2v_in0[77]),
	.c2v_77_out1(c2v_in1[77]),
	.c2v_77_out2(c2v_in2[77]),
	.c2v_77_out3(c2v_in3[77]),
	.c2v_77_out4(c2v_in4[77]),
	.c2v_77_out5(c2v_in5[77]),
	.c2v_78_out0(c2v_in0[78]),
	.c2v_78_out1(c2v_in1[78]),
	.c2v_78_out2(c2v_in2[78]),
	.c2v_78_out3(c2v_in3[78]),
	.c2v_78_out4(c2v_in4[78]),
	.c2v_78_out5(c2v_in5[78]),
	.c2v_79_out0(c2v_in0[79]),
	.c2v_79_out1(c2v_in1[79]),
	.c2v_79_out2(c2v_in2[79]),
	.c2v_79_out3(c2v_in3[79]),
	.c2v_79_out4(c2v_in4[79]),
	.c2v_79_out5(c2v_in5[79]),
	.c2v_80_out0(c2v_in0[80]),
	.c2v_80_out1(c2v_in1[80]),
	.c2v_80_out2(c2v_in2[80]),
	.c2v_80_out3(c2v_in3[80]),
	.c2v_80_out4(c2v_in4[80]),
	.c2v_80_out5(c2v_in5[80]),
	.c2v_81_out0(c2v_in0[81]),
	.c2v_81_out1(c2v_in1[81]),
	.c2v_81_out2(c2v_in2[81]),
	.c2v_81_out3(c2v_in3[81]),
	.c2v_81_out4(c2v_in4[81]),
	.c2v_81_out5(c2v_in5[81]),
	.c2v_82_out0(c2v_in0[82]),
	.c2v_82_out1(c2v_in1[82]),
	.c2v_82_out2(c2v_in2[82]),
	.c2v_82_out3(c2v_in3[82]),
	.c2v_82_out4(c2v_in4[82]),
	.c2v_82_out5(c2v_in5[82]),
	.c2v_83_out0(c2v_in0[83]),
	.c2v_83_out1(c2v_in1[83]),
	.c2v_83_out2(c2v_in2[83]),
	.c2v_83_out3(c2v_in3[83]),
	.c2v_83_out4(c2v_in4[83]),
	.c2v_83_out5(c2v_in5[83]),
	.c2v_84_out0(c2v_in0[84]),
	.c2v_84_out1(c2v_in1[84]),
	.c2v_84_out2(c2v_in2[84]),
	.c2v_84_out3(c2v_in3[84]),
	.c2v_84_out4(c2v_in4[84]),
	.c2v_84_out5(c2v_in5[84]),
	.c2v_85_out0(c2v_in0[85]),
	.c2v_85_out1(c2v_in1[85]),
	.c2v_85_out2(c2v_in2[85]),
	.c2v_85_out3(c2v_in3[85]),
	.c2v_85_out4(c2v_in4[85]),
	.c2v_85_out5(c2v_in5[85]),
	.c2v_86_out0(c2v_in0[86]),
	.c2v_86_out1(c2v_in1[86]),
	.c2v_86_out2(c2v_in2[86]),
	.c2v_86_out3(c2v_in3[86]),
	.c2v_86_out4(c2v_in4[86]),
	.c2v_86_out5(c2v_in5[86]),
	.c2v_87_out0(c2v_in0[87]),
	.c2v_87_out1(c2v_in1[87]),
	.c2v_87_out2(c2v_in2[87]),
	.c2v_87_out3(c2v_in3[87]),
	.c2v_87_out4(c2v_in4[87]),
	.c2v_87_out5(c2v_in5[87]),
	.c2v_88_out0(c2v_in0[88]),
	.c2v_88_out1(c2v_in1[88]),
	.c2v_88_out2(c2v_in2[88]),
	.c2v_88_out3(c2v_in3[88]),
	.c2v_88_out4(c2v_in4[88]),
	.c2v_88_out5(c2v_in5[88]),
	.c2v_89_out0(c2v_in0[89]),
	.c2v_89_out1(c2v_in1[89]),
	.c2v_89_out2(c2v_in2[89]),
	.c2v_89_out3(c2v_in3[89]),
	.c2v_89_out4(c2v_in4[89]),
	.c2v_89_out5(c2v_in5[89]),
	.c2v_90_out0(c2v_in0[90]),
	.c2v_90_out1(c2v_in1[90]),
	.c2v_90_out2(c2v_in2[90]),
	.c2v_90_out3(c2v_in3[90]),
	.c2v_90_out4(c2v_in4[90]),
	.c2v_90_out5(c2v_in5[90]),
	.c2v_91_out0(c2v_in0[91]),
	.c2v_91_out1(c2v_in1[91]),
	.c2v_91_out2(c2v_in2[91]),
	.c2v_91_out3(c2v_in3[91]),
	.c2v_91_out4(c2v_in4[91]),
	.c2v_91_out5(c2v_in5[91]),
	.c2v_92_out0(c2v_in0[92]),
	.c2v_92_out1(c2v_in1[92]),
	.c2v_92_out2(c2v_in2[92]),
	.c2v_92_out3(c2v_in3[92]),
	.c2v_92_out4(c2v_in4[92]),
	.c2v_92_out5(c2v_in5[92]),
	.c2v_93_out0(c2v_in0[93]),
	.c2v_93_out1(c2v_in1[93]),
	.c2v_93_out2(c2v_in2[93]),
	.c2v_93_out3(c2v_in3[93]),
	.c2v_93_out4(c2v_in4[93]),
	.c2v_93_out5(c2v_in5[93]),
	.c2v_94_out0(c2v_in0[94]),
	.c2v_94_out1(c2v_in1[94]),
	.c2v_94_out2(c2v_in2[94]),
	.c2v_94_out3(c2v_in3[94]),
	.c2v_94_out4(c2v_in4[94]),
	.c2v_94_out5(c2v_in5[94]),
	.c2v_95_out0(c2v_in0[95]),
	.c2v_95_out1(c2v_in1[95]),
	.c2v_95_out2(c2v_in2[95]),
	.c2v_95_out3(c2v_in3[95]),
	.c2v_95_out4(c2v_in4[95]),
	.c2v_95_out5(c2v_in5[95]),
	.c2v_96_out0(c2v_in0[96]),
	.c2v_96_out1(c2v_in1[96]),
	.c2v_96_out2(c2v_in2[96]),
	.c2v_96_out3(c2v_in3[96]),
	.c2v_96_out4(c2v_in4[96]),
	.c2v_96_out5(c2v_in5[96]),
	.c2v_97_out0(c2v_in0[97]),
	.c2v_97_out1(c2v_in1[97]),
	.c2v_97_out2(c2v_in2[97]),
	.c2v_97_out3(c2v_in3[97]),
	.c2v_97_out4(c2v_in4[97]),
	.c2v_97_out5(c2v_in5[97]),
	.c2v_98_out0(c2v_in0[98]),
	.c2v_98_out1(c2v_in1[98]),
	.c2v_98_out2(c2v_in2[98]),
	.c2v_98_out3(c2v_in3[98]),
	.c2v_98_out4(c2v_in4[98]),
	.c2v_98_out5(c2v_in5[98]),
	.c2v_99_out0(c2v_in0[99]),
	.c2v_99_out1(c2v_in1[99]),
	.c2v_99_out2(c2v_in2[99]),
	.c2v_99_out3(c2v_in3[99]),
	.c2v_99_out4(c2v_in4[99]),
	.c2v_99_out5(c2v_in5[99]),
	.c2v_100_out0(c2v_in0[100]),
	.c2v_100_out1(c2v_in1[100]),
	.c2v_100_out2(c2v_in2[100]),
	.c2v_100_out3(c2v_in3[100]),
	.c2v_100_out4(c2v_in4[100]),
	.c2v_100_out5(c2v_in5[100]),
	.c2v_101_out0(c2v_in0[101]),
	.c2v_101_out1(c2v_in1[101]),
	.c2v_101_out2(c2v_in2[101]),
	.c2v_101_out3(c2v_in3[101]),
	.c2v_101_out4(c2v_in4[101]),
	.c2v_101_out5(c2v_in5[101]),

	.v2c_0_in0(v2c_out0[0]),
	.v2c_0_in1(v2c_out1[0]),
	.v2c_0_in2(v2c_out2[0]),
	.v2c_0_in3(v2c_out3[0]),
	.v2c_0_in4(v2c_out4[0]),
	.v2c_0_in5(v2c_out5[0]),
	.v2c_1_in0(v2c_out0[1]),
	.v2c_1_in1(v2c_out1[1]),
	.v2c_1_in2(v2c_out2[1]),
	.v2c_1_in3(v2c_out3[1]),
	.v2c_1_in4(v2c_out4[1]),
	.v2c_1_in5(v2c_out5[1]),
	.v2c_2_in0(v2c_out0[2]),
	.v2c_2_in1(v2c_out1[2]),
	.v2c_2_in2(v2c_out2[2]),
	.v2c_2_in3(v2c_out3[2]),
	.v2c_2_in4(v2c_out4[2]),
	.v2c_2_in5(v2c_out5[2]),
	.v2c_3_in0(v2c_out0[3]),
	.v2c_3_in1(v2c_out1[3]),
	.v2c_3_in2(v2c_out2[3]),
	.v2c_3_in3(v2c_out3[3]),
	.v2c_3_in4(v2c_out4[3]),
	.v2c_3_in5(v2c_out5[3]),
	.v2c_4_in0(v2c_out0[4]),
	.v2c_4_in1(v2c_out1[4]),
	.v2c_4_in2(v2c_out2[4]),
	.v2c_4_in3(v2c_out3[4]),
	.v2c_4_in4(v2c_out4[4]),
	.v2c_4_in5(v2c_out5[4]),
	.v2c_5_in0(v2c_out0[5]),
	.v2c_5_in1(v2c_out1[5]),
	.v2c_5_in2(v2c_out2[5]),
	.v2c_5_in3(v2c_out3[5]),
	.v2c_5_in4(v2c_out4[5]),
	.v2c_5_in5(v2c_out5[5]),
	.v2c_6_in0(v2c_out0[6]),
	.v2c_6_in1(v2c_out1[6]),
	.v2c_6_in2(v2c_out2[6]),
	.v2c_6_in3(v2c_out3[6]),
	.v2c_6_in4(v2c_out4[6]),
	.v2c_6_in5(v2c_out5[6]),
	.v2c_7_in0(v2c_out0[7]),
	.v2c_7_in1(v2c_out1[7]),
	.v2c_7_in2(v2c_out2[7]),
	.v2c_7_in3(v2c_out3[7]),
	.v2c_7_in4(v2c_out4[7]),
	.v2c_7_in5(v2c_out5[7]),
	.v2c_8_in0(v2c_out0[8]),
	.v2c_8_in1(v2c_out1[8]),
	.v2c_8_in2(v2c_out2[8]),
	.v2c_8_in3(v2c_out3[8]),
	.v2c_8_in4(v2c_out4[8]),
	.v2c_8_in5(v2c_out5[8]),
	.v2c_9_in0(v2c_out0[9]),
	.v2c_9_in1(v2c_out1[9]),
	.v2c_9_in2(v2c_out2[9]),
	.v2c_9_in3(v2c_out3[9]),
	.v2c_9_in4(v2c_out4[9]),
	.v2c_9_in5(v2c_out5[9]),
	.v2c_10_in0(v2c_out0[10]),
	.v2c_10_in1(v2c_out1[10]),
	.v2c_10_in2(v2c_out2[10]),
	.v2c_10_in3(v2c_out3[10]),
	.v2c_10_in4(v2c_out4[10]),
	.v2c_10_in5(v2c_out5[10]),
	.v2c_11_in0(v2c_out0[11]),
	.v2c_11_in1(v2c_out1[11]),
	.v2c_11_in2(v2c_out2[11]),
	.v2c_11_in3(v2c_out3[11]),
	.v2c_11_in4(v2c_out4[11]),
	.v2c_11_in5(v2c_out5[11]),
	.v2c_12_in0(v2c_out0[12]),
	.v2c_12_in1(v2c_out1[12]),
	.v2c_12_in2(v2c_out2[12]),
	.v2c_12_in3(v2c_out3[12]),
	.v2c_12_in4(v2c_out4[12]),
	.v2c_12_in5(v2c_out5[12]),
	.v2c_13_in0(v2c_out0[13]),
	.v2c_13_in1(v2c_out1[13]),
	.v2c_13_in2(v2c_out2[13]),
	.v2c_13_in3(v2c_out3[13]),
	.v2c_13_in4(v2c_out4[13]),
	.v2c_13_in5(v2c_out5[13]),
	.v2c_14_in0(v2c_out0[14]),
	.v2c_14_in1(v2c_out1[14]),
	.v2c_14_in2(v2c_out2[14]),
	.v2c_14_in3(v2c_out3[14]),
	.v2c_14_in4(v2c_out4[14]),
	.v2c_14_in5(v2c_out5[14]),
	.v2c_15_in0(v2c_out0[15]),
	.v2c_15_in1(v2c_out1[15]),
	.v2c_15_in2(v2c_out2[15]),
	.v2c_15_in3(v2c_out3[15]),
	.v2c_15_in4(v2c_out4[15]),
	.v2c_15_in5(v2c_out5[15]),
	.v2c_16_in0(v2c_out0[16]),
	.v2c_16_in1(v2c_out1[16]),
	.v2c_16_in2(v2c_out2[16]),
	.v2c_16_in3(v2c_out3[16]),
	.v2c_16_in4(v2c_out4[16]),
	.v2c_16_in5(v2c_out5[16]),
	.v2c_17_in0(v2c_out0[17]),
	.v2c_17_in1(v2c_out1[17]),
	.v2c_17_in2(v2c_out2[17]),
	.v2c_17_in3(v2c_out3[17]),
	.v2c_17_in4(v2c_out4[17]),
	.v2c_17_in5(v2c_out5[17]),
	.v2c_18_in0(v2c_out0[18]),
	.v2c_18_in1(v2c_out1[18]),
	.v2c_18_in2(v2c_out2[18]),
	.v2c_18_in3(v2c_out3[18]),
	.v2c_18_in4(v2c_out4[18]),
	.v2c_18_in5(v2c_out5[18]),
	.v2c_19_in0(v2c_out0[19]),
	.v2c_19_in1(v2c_out1[19]),
	.v2c_19_in2(v2c_out2[19]),
	.v2c_19_in3(v2c_out3[19]),
	.v2c_19_in4(v2c_out4[19]),
	.v2c_19_in5(v2c_out5[19]),
	.v2c_20_in0(v2c_out0[20]),
	.v2c_20_in1(v2c_out1[20]),
	.v2c_20_in2(v2c_out2[20]),
	.v2c_20_in3(v2c_out3[20]),
	.v2c_20_in4(v2c_out4[20]),
	.v2c_20_in5(v2c_out5[20]),
	.v2c_21_in0(v2c_out0[21]),
	.v2c_21_in1(v2c_out1[21]),
	.v2c_21_in2(v2c_out2[21]),
	.v2c_21_in3(v2c_out3[21]),
	.v2c_21_in4(v2c_out4[21]),
	.v2c_21_in5(v2c_out5[21]),
	.v2c_22_in0(v2c_out0[22]),
	.v2c_22_in1(v2c_out1[22]),
	.v2c_22_in2(v2c_out2[22]),
	.v2c_22_in3(v2c_out3[22]),
	.v2c_22_in4(v2c_out4[22]),
	.v2c_22_in5(v2c_out5[22]),
	.v2c_23_in0(v2c_out0[23]),
	.v2c_23_in1(v2c_out1[23]),
	.v2c_23_in2(v2c_out2[23]),
	.v2c_23_in3(v2c_out3[23]),
	.v2c_23_in4(v2c_out4[23]),
	.v2c_23_in5(v2c_out5[23]),
	.v2c_24_in0(v2c_out0[24]),
	.v2c_24_in1(v2c_out1[24]),
	.v2c_24_in2(v2c_out2[24]),
	.v2c_24_in3(v2c_out3[24]),
	.v2c_24_in4(v2c_out4[24]),
	.v2c_24_in5(v2c_out5[24]),
	.v2c_25_in0(v2c_out0[25]),
	.v2c_25_in1(v2c_out1[25]),
	.v2c_25_in2(v2c_out2[25]),
	.v2c_25_in3(v2c_out3[25]),
	.v2c_25_in4(v2c_out4[25]),
	.v2c_25_in5(v2c_out5[25]),
	.v2c_26_in0(v2c_out0[26]),
	.v2c_26_in1(v2c_out1[26]),
	.v2c_26_in2(v2c_out2[26]),
	.v2c_26_in3(v2c_out3[26]),
	.v2c_26_in4(v2c_out4[26]),
	.v2c_26_in5(v2c_out5[26]),
	.v2c_27_in0(v2c_out0[27]),
	.v2c_27_in1(v2c_out1[27]),
	.v2c_27_in2(v2c_out2[27]),
	.v2c_27_in3(v2c_out3[27]),
	.v2c_27_in4(v2c_out4[27]),
	.v2c_27_in5(v2c_out5[27]),
	.v2c_28_in0(v2c_out0[28]),
	.v2c_28_in1(v2c_out1[28]),
	.v2c_28_in2(v2c_out2[28]),
	.v2c_28_in3(v2c_out3[28]),
	.v2c_28_in4(v2c_out4[28]),
	.v2c_28_in5(v2c_out5[28]),
	.v2c_29_in0(v2c_out0[29]),
	.v2c_29_in1(v2c_out1[29]),
	.v2c_29_in2(v2c_out2[29]),
	.v2c_29_in3(v2c_out3[29]),
	.v2c_29_in4(v2c_out4[29]),
	.v2c_29_in5(v2c_out5[29]),
	.v2c_30_in0(v2c_out0[30]),
	.v2c_30_in1(v2c_out1[30]),
	.v2c_30_in2(v2c_out2[30]),
	.v2c_30_in3(v2c_out3[30]),
	.v2c_30_in4(v2c_out4[30]),
	.v2c_30_in5(v2c_out5[30]),
	.v2c_31_in0(v2c_out0[31]),
	.v2c_31_in1(v2c_out1[31]),
	.v2c_31_in2(v2c_out2[31]),
	.v2c_31_in3(v2c_out3[31]),
	.v2c_31_in4(v2c_out4[31]),
	.v2c_31_in5(v2c_out5[31]),
	.v2c_32_in0(v2c_out0[32]),
	.v2c_32_in1(v2c_out1[32]),
	.v2c_32_in2(v2c_out2[32]),
	.v2c_32_in3(v2c_out3[32]),
	.v2c_32_in4(v2c_out4[32]),
	.v2c_32_in5(v2c_out5[32]),
	.v2c_33_in0(v2c_out0[33]),
	.v2c_33_in1(v2c_out1[33]),
	.v2c_33_in2(v2c_out2[33]),
	.v2c_33_in3(v2c_out3[33]),
	.v2c_33_in4(v2c_out4[33]),
	.v2c_33_in5(v2c_out5[33]),
	.v2c_34_in0(v2c_out0[34]),
	.v2c_34_in1(v2c_out1[34]),
	.v2c_34_in2(v2c_out2[34]),
	.v2c_34_in3(v2c_out3[34]),
	.v2c_34_in4(v2c_out4[34]),
	.v2c_34_in5(v2c_out5[34]),
	.v2c_35_in0(v2c_out0[35]),
	.v2c_35_in1(v2c_out1[35]),
	.v2c_35_in2(v2c_out2[35]),
	.v2c_35_in3(v2c_out3[35]),
	.v2c_35_in4(v2c_out4[35]),
	.v2c_35_in5(v2c_out5[35]),
	.v2c_36_in0(v2c_out0[36]),
	.v2c_36_in1(v2c_out1[36]),
	.v2c_36_in2(v2c_out2[36]),
	.v2c_36_in3(v2c_out3[36]),
	.v2c_36_in4(v2c_out4[36]),
	.v2c_36_in5(v2c_out5[36]),
	.v2c_37_in0(v2c_out0[37]),
	.v2c_37_in1(v2c_out1[37]),
	.v2c_37_in2(v2c_out2[37]),
	.v2c_37_in3(v2c_out3[37]),
	.v2c_37_in4(v2c_out4[37]),
	.v2c_37_in5(v2c_out5[37]),
	.v2c_38_in0(v2c_out0[38]),
	.v2c_38_in1(v2c_out1[38]),
	.v2c_38_in2(v2c_out2[38]),
	.v2c_38_in3(v2c_out3[38]),
	.v2c_38_in4(v2c_out4[38]),
	.v2c_38_in5(v2c_out5[38]),
	.v2c_39_in0(v2c_out0[39]),
	.v2c_39_in1(v2c_out1[39]),
	.v2c_39_in2(v2c_out2[39]),
	.v2c_39_in3(v2c_out3[39]),
	.v2c_39_in4(v2c_out4[39]),
	.v2c_39_in5(v2c_out5[39]),
	.v2c_40_in0(v2c_out0[40]),
	.v2c_40_in1(v2c_out1[40]),
	.v2c_40_in2(v2c_out2[40]),
	.v2c_40_in3(v2c_out3[40]),
	.v2c_40_in4(v2c_out4[40]),
	.v2c_40_in5(v2c_out5[40]),
	.v2c_41_in0(v2c_out0[41]),
	.v2c_41_in1(v2c_out1[41]),
	.v2c_41_in2(v2c_out2[41]),
	.v2c_41_in3(v2c_out3[41]),
	.v2c_41_in4(v2c_out4[41]),
	.v2c_41_in5(v2c_out5[41]),
	.v2c_42_in0(v2c_out0[42]),
	.v2c_42_in1(v2c_out1[42]),
	.v2c_42_in2(v2c_out2[42]),
	.v2c_42_in3(v2c_out3[42]),
	.v2c_42_in4(v2c_out4[42]),
	.v2c_42_in5(v2c_out5[42]),
	.v2c_43_in0(v2c_out0[43]),
	.v2c_43_in1(v2c_out1[43]),
	.v2c_43_in2(v2c_out2[43]),
	.v2c_43_in3(v2c_out3[43]),
	.v2c_43_in4(v2c_out4[43]),
	.v2c_43_in5(v2c_out5[43]),
	.v2c_44_in0(v2c_out0[44]),
	.v2c_44_in1(v2c_out1[44]),
	.v2c_44_in2(v2c_out2[44]),
	.v2c_44_in3(v2c_out3[44]),
	.v2c_44_in4(v2c_out4[44]),
	.v2c_44_in5(v2c_out5[44]),
	.v2c_45_in0(v2c_out0[45]),
	.v2c_45_in1(v2c_out1[45]),
	.v2c_45_in2(v2c_out2[45]),
	.v2c_45_in3(v2c_out3[45]),
	.v2c_45_in4(v2c_out4[45]),
	.v2c_45_in5(v2c_out5[45]),
	.v2c_46_in0(v2c_out0[46]),
	.v2c_46_in1(v2c_out1[46]),
	.v2c_46_in2(v2c_out2[46]),
	.v2c_46_in3(v2c_out3[46]),
	.v2c_46_in4(v2c_out4[46]),
	.v2c_46_in5(v2c_out5[46]),
	.v2c_47_in0(v2c_out0[47]),
	.v2c_47_in1(v2c_out1[47]),
	.v2c_47_in2(v2c_out2[47]),
	.v2c_47_in3(v2c_out3[47]),
	.v2c_47_in4(v2c_out4[47]),
	.v2c_47_in5(v2c_out5[47]),
	.v2c_48_in0(v2c_out0[48]),
	.v2c_48_in1(v2c_out1[48]),
	.v2c_48_in2(v2c_out2[48]),
	.v2c_48_in3(v2c_out3[48]),
	.v2c_48_in4(v2c_out4[48]),
	.v2c_48_in5(v2c_out5[48]),
	.v2c_49_in0(v2c_out0[49]),
	.v2c_49_in1(v2c_out1[49]),
	.v2c_49_in2(v2c_out2[49]),
	.v2c_49_in3(v2c_out3[49]),
	.v2c_49_in4(v2c_out4[49]),
	.v2c_49_in5(v2c_out5[49]),
	.v2c_50_in0(v2c_out0[50]),
	.v2c_50_in1(v2c_out1[50]),
	.v2c_50_in2(v2c_out2[50]),
	.v2c_50_in3(v2c_out3[50]),
	.v2c_50_in4(v2c_out4[50]),
	.v2c_50_in5(v2c_out5[50]),
	.v2c_51_in0(v2c_out0[51]),
	.v2c_51_in1(v2c_out1[51]),
	.v2c_51_in2(v2c_out2[51]),
	.v2c_51_in3(v2c_out3[51]),
	.v2c_51_in4(v2c_out4[51]),
	.v2c_51_in5(v2c_out5[51]),
	.v2c_52_in0(v2c_out0[52]),
	.v2c_52_in1(v2c_out1[52]),
	.v2c_52_in2(v2c_out2[52]),
	.v2c_52_in3(v2c_out3[52]),
	.v2c_52_in4(v2c_out4[52]),
	.v2c_52_in5(v2c_out5[52]),
	.v2c_53_in0(v2c_out0[53]),
	.v2c_53_in1(v2c_out1[53]),
	.v2c_53_in2(v2c_out2[53]),
	.v2c_53_in3(v2c_out3[53]),
	.v2c_53_in4(v2c_out4[53]),
	.v2c_53_in5(v2c_out5[53]),
	.v2c_54_in0(v2c_out0[54]),
	.v2c_54_in1(v2c_out1[54]),
	.v2c_54_in2(v2c_out2[54]),
	.v2c_54_in3(v2c_out3[54]),
	.v2c_54_in4(v2c_out4[54]),
	.v2c_54_in5(v2c_out5[54]),
	.v2c_55_in0(v2c_out0[55]),
	.v2c_55_in1(v2c_out1[55]),
	.v2c_55_in2(v2c_out2[55]),
	.v2c_55_in3(v2c_out3[55]),
	.v2c_55_in4(v2c_out4[55]),
	.v2c_55_in5(v2c_out5[55]),
	.v2c_56_in0(v2c_out0[56]),
	.v2c_56_in1(v2c_out1[56]),
	.v2c_56_in2(v2c_out2[56]),
	.v2c_56_in3(v2c_out3[56]),
	.v2c_56_in4(v2c_out4[56]),
	.v2c_56_in5(v2c_out5[56]),
	.v2c_57_in0(v2c_out0[57]),
	.v2c_57_in1(v2c_out1[57]),
	.v2c_57_in2(v2c_out2[57]),
	.v2c_57_in3(v2c_out3[57]),
	.v2c_57_in4(v2c_out4[57]),
	.v2c_57_in5(v2c_out5[57]),
	.v2c_58_in0(v2c_out0[58]),
	.v2c_58_in1(v2c_out1[58]),
	.v2c_58_in2(v2c_out2[58]),
	.v2c_58_in3(v2c_out3[58]),
	.v2c_58_in4(v2c_out4[58]),
	.v2c_58_in5(v2c_out5[58]),
	.v2c_59_in0(v2c_out0[59]),
	.v2c_59_in1(v2c_out1[59]),
	.v2c_59_in2(v2c_out2[59]),
	.v2c_59_in3(v2c_out3[59]),
	.v2c_59_in4(v2c_out4[59]),
	.v2c_59_in5(v2c_out5[59]),
	.v2c_60_in0(v2c_out0[60]),
	.v2c_60_in1(v2c_out1[60]),
	.v2c_60_in2(v2c_out2[60]),
	.v2c_60_in3(v2c_out3[60]),
	.v2c_60_in4(v2c_out4[60]),
	.v2c_60_in5(v2c_out5[60]),
	.v2c_61_in0(v2c_out0[61]),
	.v2c_61_in1(v2c_out1[61]),
	.v2c_61_in2(v2c_out2[61]),
	.v2c_61_in3(v2c_out3[61]),
	.v2c_61_in4(v2c_out4[61]),
	.v2c_61_in5(v2c_out5[61]),
	.v2c_62_in0(v2c_out0[62]),
	.v2c_62_in1(v2c_out1[62]),
	.v2c_62_in2(v2c_out2[62]),
	.v2c_62_in3(v2c_out3[62]),
	.v2c_62_in4(v2c_out4[62]),
	.v2c_62_in5(v2c_out5[62]),
	.v2c_63_in0(v2c_out0[63]),
	.v2c_63_in1(v2c_out1[63]),
	.v2c_63_in2(v2c_out2[63]),
	.v2c_63_in3(v2c_out3[63]),
	.v2c_63_in4(v2c_out4[63]),
	.v2c_63_in5(v2c_out5[63]),
	.v2c_64_in0(v2c_out0[64]),
	.v2c_64_in1(v2c_out1[64]),
	.v2c_64_in2(v2c_out2[64]),
	.v2c_64_in3(v2c_out3[64]),
	.v2c_64_in4(v2c_out4[64]),
	.v2c_64_in5(v2c_out5[64]),
	.v2c_65_in0(v2c_out0[65]),
	.v2c_65_in1(v2c_out1[65]),
	.v2c_65_in2(v2c_out2[65]),
	.v2c_65_in3(v2c_out3[65]),
	.v2c_65_in4(v2c_out4[65]),
	.v2c_65_in5(v2c_out5[65]),
	.v2c_66_in0(v2c_out0[66]),
	.v2c_66_in1(v2c_out1[66]),
	.v2c_66_in2(v2c_out2[66]),
	.v2c_66_in3(v2c_out3[66]),
	.v2c_66_in4(v2c_out4[66]),
	.v2c_66_in5(v2c_out5[66]),
	.v2c_67_in0(v2c_out0[67]),
	.v2c_67_in1(v2c_out1[67]),
	.v2c_67_in2(v2c_out2[67]),
	.v2c_67_in3(v2c_out3[67]),
	.v2c_67_in4(v2c_out4[67]),
	.v2c_67_in5(v2c_out5[67]),
	.v2c_68_in0(v2c_out0[68]),
	.v2c_68_in1(v2c_out1[68]),
	.v2c_68_in2(v2c_out2[68]),
	.v2c_68_in3(v2c_out3[68]),
	.v2c_68_in4(v2c_out4[68]),
	.v2c_68_in5(v2c_out5[68]),
	.v2c_69_in0(v2c_out0[69]),
	.v2c_69_in1(v2c_out1[69]),
	.v2c_69_in2(v2c_out2[69]),
	.v2c_69_in3(v2c_out3[69]),
	.v2c_69_in4(v2c_out4[69]),
	.v2c_69_in5(v2c_out5[69]),
	.v2c_70_in0(v2c_out0[70]),
	.v2c_70_in1(v2c_out1[70]),
	.v2c_70_in2(v2c_out2[70]),
	.v2c_70_in3(v2c_out3[70]),
	.v2c_70_in4(v2c_out4[70]),
	.v2c_70_in5(v2c_out5[70]),
	.v2c_71_in0(v2c_out0[71]),
	.v2c_71_in1(v2c_out1[71]),
	.v2c_71_in2(v2c_out2[71]),
	.v2c_71_in3(v2c_out3[71]),
	.v2c_71_in4(v2c_out4[71]),
	.v2c_71_in5(v2c_out5[71]),
	.v2c_72_in0(v2c_out0[72]),
	.v2c_72_in1(v2c_out1[72]),
	.v2c_72_in2(v2c_out2[72]),
	.v2c_72_in3(v2c_out3[72]),
	.v2c_72_in4(v2c_out4[72]),
	.v2c_72_in5(v2c_out5[72]),
	.v2c_73_in0(v2c_out0[73]),
	.v2c_73_in1(v2c_out1[73]),
	.v2c_73_in2(v2c_out2[73]),
	.v2c_73_in3(v2c_out3[73]),
	.v2c_73_in4(v2c_out4[73]),
	.v2c_73_in5(v2c_out5[73]),
	.v2c_74_in0(v2c_out0[74]),
	.v2c_74_in1(v2c_out1[74]),
	.v2c_74_in2(v2c_out2[74]),
	.v2c_74_in3(v2c_out3[74]),
	.v2c_74_in4(v2c_out4[74]),
	.v2c_74_in5(v2c_out5[74]),
	.v2c_75_in0(v2c_out0[75]),
	.v2c_75_in1(v2c_out1[75]),
	.v2c_75_in2(v2c_out2[75]),
	.v2c_75_in3(v2c_out3[75]),
	.v2c_75_in4(v2c_out4[75]),
	.v2c_75_in5(v2c_out5[75]),
	.v2c_76_in0(v2c_out0[76]),
	.v2c_76_in1(v2c_out1[76]),
	.v2c_76_in2(v2c_out2[76]),
	.v2c_76_in3(v2c_out3[76]),
	.v2c_76_in4(v2c_out4[76]),
	.v2c_76_in5(v2c_out5[76]),
	.v2c_77_in0(v2c_out0[77]),
	.v2c_77_in1(v2c_out1[77]),
	.v2c_77_in2(v2c_out2[77]),
	.v2c_77_in3(v2c_out3[77]),
	.v2c_77_in4(v2c_out4[77]),
	.v2c_77_in5(v2c_out5[77]),
	.v2c_78_in0(v2c_out0[78]),
	.v2c_78_in1(v2c_out1[78]),
	.v2c_78_in2(v2c_out2[78]),
	.v2c_78_in3(v2c_out3[78]),
	.v2c_78_in4(v2c_out4[78]),
	.v2c_78_in5(v2c_out5[78]),
	.v2c_79_in0(v2c_out0[79]),
	.v2c_79_in1(v2c_out1[79]),
	.v2c_79_in2(v2c_out2[79]),
	.v2c_79_in3(v2c_out3[79]),
	.v2c_79_in4(v2c_out4[79]),
	.v2c_79_in5(v2c_out5[79]),
	.v2c_80_in0(v2c_out0[80]),
	.v2c_80_in1(v2c_out1[80]),
	.v2c_80_in2(v2c_out2[80]),
	.v2c_80_in3(v2c_out3[80]),
	.v2c_80_in4(v2c_out4[80]),
	.v2c_80_in5(v2c_out5[80]),
	.v2c_81_in0(v2c_out0[81]),
	.v2c_81_in1(v2c_out1[81]),
	.v2c_81_in2(v2c_out2[81]),
	.v2c_81_in3(v2c_out3[81]),
	.v2c_81_in4(v2c_out4[81]),
	.v2c_81_in5(v2c_out5[81]),
	.v2c_82_in0(v2c_out0[82]),
	.v2c_82_in1(v2c_out1[82]),
	.v2c_82_in2(v2c_out2[82]),
	.v2c_82_in3(v2c_out3[82]),
	.v2c_82_in4(v2c_out4[82]),
	.v2c_82_in5(v2c_out5[82]),
	.v2c_83_in0(v2c_out0[83]),
	.v2c_83_in1(v2c_out1[83]),
	.v2c_83_in2(v2c_out2[83]),
	.v2c_83_in3(v2c_out3[83]),
	.v2c_83_in4(v2c_out4[83]),
	.v2c_83_in5(v2c_out5[83]),
	.v2c_84_in0(v2c_out0[84]),
	.v2c_84_in1(v2c_out1[84]),
	.v2c_84_in2(v2c_out2[84]),
	.v2c_84_in3(v2c_out3[84]),
	.v2c_84_in4(v2c_out4[84]),
	.v2c_84_in5(v2c_out5[84]),
	.v2c_85_in0(v2c_out0[85]),
	.v2c_85_in1(v2c_out1[85]),
	.v2c_85_in2(v2c_out2[85]),
	.v2c_85_in3(v2c_out3[85]),
	.v2c_85_in4(v2c_out4[85]),
	.v2c_85_in5(v2c_out5[85]),
	.v2c_86_in0(v2c_out0[86]),
	.v2c_86_in1(v2c_out1[86]),
	.v2c_86_in2(v2c_out2[86]),
	.v2c_86_in3(v2c_out3[86]),
	.v2c_86_in4(v2c_out4[86]),
	.v2c_86_in5(v2c_out5[86]),
	.v2c_87_in0(v2c_out0[87]),
	.v2c_87_in1(v2c_out1[87]),
	.v2c_87_in2(v2c_out2[87]),
	.v2c_87_in3(v2c_out3[87]),
	.v2c_87_in4(v2c_out4[87]),
	.v2c_87_in5(v2c_out5[87]),
	.v2c_88_in0(v2c_out0[88]),
	.v2c_88_in1(v2c_out1[88]),
	.v2c_88_in2(v2c_out2[88]),
	.v2c_88_in3(v2c_out3[88]),
	.v2c_88_in4(v2c_out4[88]),
	.v2c_88_in5(v2c_out5[88]),
	.v2c_89_in0(v2c_out0[89]),
	.v2c_89_in1(v2c_out1[89]),
	.v2c_89_in2(v2c_out2[89]),
	.v2c_89_in3(v2c_out3[89]),
	.v2c_89_in4(v2c_out4[89]),
	.v2c_89_in5(v2c_out5[89]),
	.v2c_90_in0(v2c_out0[90]),
	.v2c_90_in1(v2c_out1[90]),
	.v2c_90_in2(v2c_out2[90]),
	.v2c_90_in3(v2c_out3[90]),
	.v2c_90_in4(v2c_out4[90]),
	.v2c_90_in5(v2c_out5[90]),
	.v2c_91_in0(v2c_out0[91]),
	.v2c_91_in1(v2c_out1[91]),
	.v2c_91_in2(v2c_out2[91]),
	.v2c_91_in3(v2c_out3[91]),
	.v2c_91_in4(v2c_out4[91]),
	.v2c_91_in5(v2c_out5[91]),
	.v2c_92_in0(v2c_out0[92]),
	.v2c_92_in1(v2c_out1[92]),
	.v2c_92_in2(v2c_out2[92]),
	.v2c_92_in3(v2c_out3[92]),
	.v2c_92_in4(v2c_out4[92]),
	.v2c_92_in5(v2c_out5[92]),
	.v2c_93_in0(v2c_out0[93]),
	.v2c_93_in1(v2c_out1[93]),
	.v2c_93_in2(v2c_out2[93]),
	.v2c_93_in3(v2c_out3[93]),
	.v2c_93_in4(v2c_out4[93]),
	.v2c_93_in5(v2c_out5[93]),
	.v2c_94_in0(v2c_out0[94]),
	.v2c_94_in1(v2c_out1[94]),
	.v2c_94_in2(v2c_out2[94]),
	.v2c_94_in3(v2c_out3[94]),
	.v2c_94_in4(v2c_out4[94]),
	.v2c_94_in5(v2c_out5[94]),
	.v2c_95_in0(v2c_out0[95]),
	.v2c_95_in1(v2c_out1[95]),
	.v2c_95_in2(v2c_out2[95]),
	.v2c_95_in3(v2c_out3[95]),
	.v2c_95_in4(v2c_out4[95]),
	.v2c_95_in5(v2c_out5[95]),
	.v2c_96_in0(v2c_out0[96]),
	.v2c_96_in1(v2c_out1[96]),
	.v2c_96_in2(v2c_out2[96]),
	.v2c_96_in3(v2c_out3[96]),
	.v2c_96_in4(v2c_out4[96]),
	.v2c_96_in5(v2c_out5[96]),
	.v2c_97_in0(v2c_out0[97]),
	.v2c_97_in1(v2c_out1[97]),
	.v2c_97_in2(v2c_out2[97]),
	.v2c_97_in3(v2c_out3[97]),
	.v2c_97_in4(v2c_out4[97]),
	.v2c_97_in5(v2c_out5[97]),
	.v2c_98_in0(v2c_out0[98]),
	.v2c_98_in1(v2c_out1[98]),
	.v2c_98_in2(v2c_out2[98]),
	.v2c_98_in3(v2c_out3[98]),
	.v2c_98_in4(v2c_out4[98]),
	.v2c_98_in5(v2c_out5[98]),
	.v2c_99_in0(v2c_out0[99]),
	.v2c_99_in1(v2c_out1[99]),
	.v2c_99_in2(v2c_out2[99]),
	.v2c_99_in3(v2c_out3[99]),
	.v2c_99_in4(v2c_out4[99]),
	.v2c_99_in5(v2c_out5[99]),
	.v2c_100_in0(v2c_out0[100]),
	.v2c_100_in1(v2c_out1[100]),
	.v2c_100_in2(v2c_out2[100]),
	.v2c_100_in3(v2c_out3[100]),
	.v2c_100_in4(v2c_out4[100]),
	.v2c_100_in5(v2c_out5[100]),
	.v2c_101_in0(v2c_out0[101]),
	.v2c_101_in1(v2c_out1[101]),
	.v2c_101_in2(v2c_out2[101]),
	.v2c_101_in3(v2c_out3[101]),
	.v2c_101_in4(v2c_out4[101]),
	.v2c_101_in5(v2c_out5[101]),

	.read_clk (read_clk),
	.read_addr_offset (cnu_read_addr_offset),
	.v2c_latch_en (v2c_latch_en),
	.v2c_parallel_load (load[1]),

	// Iteration-Refresh Page Address
	.page_addr_ram_0(cnu_page_addr_ram_0[CN_PAGE_ADDR_BW+1-1:0]),
	.page_addr_ram_1(cnu_page_addr_ram_1[CN_PAGE_ADDR_BW+1-1:0]),
	.page_addr_ram_2(cnu_page_addr_ram_2[CN_PAGE_ADDR_BW+1-1:0]),
	.page_addr_ram_3(cnu_page_addr_ram_3[CN_PAGE_ADDR_BW+1-1:0]),
	//Iteration-Refresh Page Data
	. ram_write_dataA_0 (cnu_ram_write_dataA_0[CN_ROM_RD_BW-1:0]), // from portA of IB-ROM
	. ram_write_dataB_0 (cnu_ram_write_dataB_0[CN_ROM_RD_BW-1:0]), // from portB of IB-ROM
	. ram_write_dataA_1 (cnu_ram_write_dataA_1[CN_ROM_RD_BW-1:0]), // from portA of IB-ROM
	. ram_write_dataB_1 (cnu_ram_write_dataB_1[CN_ROM_RD_BW-1:0]), // from portB of IB-ROM
	. ram_write_dataA_2 (cnu_ram_write_dataA_2[CN_ROM_RD_BW-1:0]), // from portA of IB-ROM
	. ram_write_dataB_2 (cnu_ram_write_dataB_2[CN_ROM_RD_BW-1:0]), // from portB of IB-ROM
	. ram_write_dataA_3 (cnu_ram_write_dataA_3[CN_ROM_RD_BW-1:0]), // from portA of IB-ROM
	. ram_write_dataB_3 (cnu_ram_write_dataB_3[CN_ROM_RD_BW-1:0]), // from portB of IB-ROM
	.ib_ram_we (cnu_ib_ram_we[IB_CNU_DECOMP_funNum-1:0]),
	.write_clk (cn_write_clk)
);

// Instantiation of VNU IB-RAM wrapper
vnu3_ib_ram_wrapper #(
	.VN_ROM_RD_BW          (VN_ROM_RD_BW          ),
	.VN_ROM_ADDR_BW        (VN_ROM_ADDR_BW        ),
	.VN_PAGE_ADDR_BW       (VN_PAGE_ADDR_BW       ),
	.DN_ROM_RD_BW          (DN_ROM_RD_BW          ),
	.DN_ROM_ADDR_BW        (DN_ROM_ADDR_BW        ),
	.DN_PAGE_ADDR_BW       (DN_PAGE_ADDR_BW       ),
	.VN_DEGREE             (VN_DEGREE             ),
	.IB_VNU_DECOMP_funNum  (IB_VNU_DECOMP_funNum  ),
	.VN_NUM                (VN_NUM                ),
	.VNU3_INSTANTIATE_NUM  (VNU3_INSTANTIATE_NUM  ),
	.VNU3_INSTANTIATE_UNIT (VNU3_INSTANTIATE_UNIT ),
	.QUAN_SIZE             (QUAN_SIZE             ),
	.DATAPATH_WIDTH        (DATAPATH_WIDTH        )
) vnu_ib_ram_wrapper_u0(
	.hard_decision_0 (hard_decision[0]),
	.v2c_0_out0 (v2c_in0[0]),
	.v2c_0_out1 (v2c_in1[0]),
	.v2c_0_out2 (v2c_in2[0]),
	.hard_decision_1 (hard_decision[1]),
	.v2c_1_out0 (v2c_in0[1]),
	.v2c_1_out1 (v2c_in1[1]),
	.v2c_1_out2 (v2c_in2[1]),
	.hard_decision_2 (hard_decision[2]),
	.v2c_2_out0 (v2c_in0[2]),
	.v2c_2_out1 (v2c_in1[2]),
	.v2c_2_out2 (v2c_in2[2]),
	.hard_decision_3 (hard_decision[3]),
	.v2c_3_out0 (v2c_in0[3]),
	.v2c_3_out1 (v2c_in1[3]),
	.v2c_3_out2 (v2c_in2[3]),
	.hard_decision_4 (hard_decision[4]),
	.v2c_4_out0 (v2c_in0[4]),
	.v2c_4_out1 (v2c_in1[4]),
	.v2c_4_out2 (v2c_in2[4]),
	.hard_decision_5 (hard_decision[5]),
	.v2c_5_out0 (v2c_in0[5]),
	.v2c_5_out1 (v2c_in1[5]),
	.v2c_5_out2 (v2c_in2[5]),
	.hard_decision_6 (hard_decision[6]),
	.v2c_6_out0 (v2c_in0[6]),
	.v2c_6_out1 (v2c_in1[6]),
	.v2c_6_out2 (v2c_in2[6]),
	.hard_decision_7 (hard_decision[7]),
	.v2c_7_out0 (v2c_in0[7]),
	.v2c_7_out1 (v2c_in1[7]),
	.v2c_7_out2 (v2c_in2[7]),
	.hard_decision_8 (hard_decision[8]),
	.v2c_8_out0 (v2c_in0[8]),
	.v2c_8_out1 (v2c_in1[8]),
	.v2c_8_out2 (v2c_in2[8]),
	.hard_decision_9 (hard_decision[9]),
	.v2c_9_out0 (v2c_in0[9]),
	.v2c_9_out1 (v2c_in1[9]),
	.v2c_9_out2 (v2c_in2[9]),
	.hard_decision_10 (hard_decision[10]),
	.v2c_10_out0 (v2c_in0[10]),
	.v2c_10_out1 (v2c_in1[10]),
	.v2c_10_out2 (v2c_in2[10]),
	.hard_decision_11 (hard_decision[11]),
	.v2c_11_out0 (v2c_in0[11]),
	.v2c_11_out1 (v2c_in1[11]),
	.v2c_11_out2 (v2c_in2[11]),
	.hard_decision_12 (hard_decision[12]),
	.v2c_12_out0 (v2c_in0[12]),
	.v2c_12_out1 (v2c_in1[12]),
	.v2c_12_out2 (v2c_in2[12]),
	.hard_decision_13 (hard_decision[13]),
	.v2c_13_out0 (v2c_in0[13]),
	.v2c_13_out1 (v2c_in1[13]),
	.v2c_13_out2 (v2c_in2[13]),
	.hard_decision_14 (hard_decision[14]),
	.v2c_14_out0 (v2c_in0[14]),
	.v2c_14_out1 (v2c_in1[14]),
	.v2c_14_out2 (v2c_in2[14]),
	.hard_decision_15 (hard_decision[15]),
	.v2c_15_out0 (v2c_in0[15]),
	.v2c_15_out1 (v2c_in1[15]),
	.v2c_15_out2 (v2c_in2[15]),
	.hard_decision_16 (hard_decision[16]),
	.v2c_16_out0 (v2c_in0[16]),
	.v2c_16_out1 (v2c_in1[16]),
	.v2c_16_out2 (v2c_in2[16]),
	.hard_decision_17 (hard_decision[17]),
	.v2c_17_out0 (v2c_in0[17]),
	.v2c_17_out1 (v2c_in1[17]),
	.v2c_17_out2 (v2c_in2[17]),
	.hard_decision_18 (hard_decision[18]),
	.v2c_18_out0 (v2c_in0[18]),
	.v2c_18_out1 (v2c_in1[18]),
	.v2c_18_out2 (v2c_in2[18]),
	.hard_decision_19 (hard_decision[19]),
	.v2c_19_out0 (v2c_in0[19]),
	.v2c_19_out1 (v2c_in1[19]),
	.v2c_19_out2 (v2c_in2[19]),
	.hard_decision_20 (hard_decision[20]),
	.v2c_20_out0 (v2c_in0[20]),
	.v2c_20_out1 (v2c_in1[20]),
	.v2c_20_out2 (v2c_in2[20]),
	.hard_decision_21 (hard_decision[21]),
	.v2c_21_out0 (v2c_in0[21]),
	.v2c_21_out1 (v2c_in1[21]),
	.v2c_21_out2 (v2c_in2[21]),
	.hard_decision_22 (hard_decision[22]),
	.v2c_22_out0 (v2c_in0[22]),
	.v2c_22_out1 (v2c_in1[22]),
	.v2c_22_out2 (v2c_in2[22]),
	.hard_decision_23 (hard_decision[23]),
	.v2c_23_out0 (v2c_in0[23]),
	.v2c_23_out1 (v2c_in1[23]),
	.v2c_23_out2 (v2c_in2[23]),
	.hard_decision_24 (hard_decision[24]),
	.v2c_24_out0 (v2c_in0[24]),
	.v2c_24_out1 (v2c_in1[24]),
	.v2c_24_out2 (v2c_in2[24]),
	.hard_decision_25 (hard_decision[25]),
	.v2c_25_out0 (v2c_in0[25]),
	.v2c_25_out1 (v2c_in1[25]),
	.v2c_25_out2 (v2c_in2[25]),
	.hard_decision_26 (hard_decision[26]),
	.v2c_26_out0 (v2c_in0[26]),
	.v2c_26_out1 (v2c_in1[26]),
	.v2c_26_out2 (v2c_in2[26]),
	.hard_decision_27 (hard_decision[27]),
	.v2c_27_out0 (v2c_in0[27]),
	.v2c_27_out1 (v2c_in1[27]),
	.v2c_27_out2 (v2c_in2[27]),
	.hard_decision_28 (hard_decision[28]),
	.v2c_28_out0 (v2c_in0[28]),
	.v2c_28_out1 (v2c_in1[28]),
	.v2c_28_out2 (v2c_in2[28]),
	.hard_decision_29 (hard_decision[29]),
	.v2c_29_out0 (v2c_in0[29]),
	.v2c_29_out1 (v2c_in1[29]),
	.v2c_29_out2 (v2c_in2[29]),
	.hard_decision_30 (hard_decision[30]),
	.v2c_30_out0 (v2c_in0[30]),
	.v2c_30_out1 (v2c_in1[30]),
	.v2c_30_out2 (v2c_in2[30]),
	.hard_decision_31 (hard_decision[31]),
	.v2c_31_out0 (v2c_in0[31]),
	.v2c_31_out1 (v2c_in1[31]),
	.v2c_31_out2 (v2c_in2[31]),
	.hard_decision_32 (hard_decision[32]),
	.v2c_32_out0 (v2c_in0[32]),
	.v2c_32_out1 (v2c_in1[32]),
	.v2c_32_out2 (v2c_in2[32]),
	.hard_decision_33 (hard_decision[33]),
	.v2c_33_out0 (v2c_in0[33]),
	.v2c_33_out1 (v2c_in1[33]),
	.v2c_33_out2 (v2c_in2[33]),
	.hard_decision_34 (hard_decision[34]),
	.v2c_34_out0 (v2c_in0[34]),
	.v2c_34_out1 (v2c_in1[34]),
	.v2c_34_out2 (v2c_in2[34]),
	.hard_decision_35 (hard_decision[35]),
	.v2c_35_out0 (v2c_in0[35]),
	.v2c_35_out1 (v2c_in1[35]),
	.v2c_35_out2 (v2c_in2[35]),
	.hard_decision_36 (hard_decision[36]),
	.v2c_36_out0 (v2c_in0[36]),
	.v2c_36_out1 (v2c_in1[36]),
	.v2c_36_out2 (v2c_in2[36]),
	.hard_decision_37 (hard_decision[37]),
	.v2c_37_out0 (v2c_in0[37]),
	.v2c_37_out1 (v2c_in1[37]),
	.v2c_37_out2 (v2c_in2[37]),
	.hard_decision_38 (hard_decision[38]),
	.v2c_38_out0 (v2c_in0[38]),
	.v2c_38_out1 (v2c_in1[38]),
	.v2c_38_out2 (v2c_in2[38]),
	.hard_decision_39 (hard_decision[39]),
	.v2c_39_out0 (v2c_in0[39]),
	.v2c_39_out1 (v2c_in1[39]),
	.v2c_39_out2 (v2c_in2[39]),
	.hard_decision_40 (hard_decision[40]),
	.v2c_40_out0 (v2c_in0[40]),
	.v2c_40_out1 (v2c_in1[40]),
	.v2c_40_out2 (v2c_in2[40]),
	.hard_decision_41 (hard_decision[41]),
	.v2c_41_out0 (v2c_in0[41]),
	.v2c_41_out1 (v2c_in1[41]),
	.v2c_41_out2 (v2c_in2[41]),
	.hard_decision_42 (hard_decision[42]),
	.v2c_42_out0 (v2c_in0[42]),
	.v2c_42_out1 (v2c_in1[42]),
	.v2c_42_out2 (v2c_in2[42]),
	.hard_decision_43 (hard_decision[43]),
	.v2c_43_out0 (v2c_in0[43]),
	.v2c_43_out1 (v2c_in1[43]),
	.v2c_43_out2 (v2c_in2[43]),
	.hard_decision_44 (hard_decision[44]),
	.v2c_44_out0 (v2c_in0[44]),
	.v2c_44_out1 (v2c_in1[44]),
	.v2c_44_out2 (v2c_in2[44]),
	.hard_decision_45 (hard_decision[45]),
	.v2c_45_out0 (v2c_in0[45]),
	.v2c_45_out1 (v2c_in1[45]),
	.v2c_45_out2 (v2c_in2[45]),
	.hard_decision_46 (hard_decision[46]),
	.v2c_46_out0 (v2c_in0[46]),
	.v2c_46_out1 (v2c_in1[46]),
	.v2c_46_out2 (v2c_in2[46]),
	.hard_decision_47 (hard_decision[47]),
	.v2c_47_out0 (v2c_in0[47]),
	.v2c_47_out1 (v2c_in1[47]),
	.v2c_47_out2 (v2c_in2[47]),
	.hard_decision_48 (hard_decision[48]),
	.v2c_48_out0 (v2c_in0[48]),
	.v2c_48_out1 (v2c_in1[48]),
	.v2c_48_out2 (v2c_in2[48]),
	.hard_decision_49 (hard_decision[49]),
	.v2c_49_out0 (v2c_in0[49]),
	.v2c_49_out1 (v2c_in1[49]),
	.v2c_49_out2 (v2c_in2[49]),
	.hard_decision_50 (hard_decision[50]),
	.v2c_50_out0 (v2c_in0[50]),
	.v2c_50_out1 (v2c_in1[50]),
	.v2c_50_out2 (v2c_in2[50]),
	.hard_decision_51 (hard_decision[51]),
	.v2c_51_out0 (v2c_in0[51]),
	.v2c_51_out1 (v2c_in1[51]),
	.v2c_51_out2 (v2c_in2[51]),
	.hard_decision_52 (hard_decision[52]),
	.v2c_52_out0 (v2c_in0[52]),
	.v2c_52_out1 (v2c_in1[52]),
	.v2c_52_out2 (v2c_in2[52]),
	.hard_decision_53 (hard_decision[53]),
	.v2c_53_out0 (v2c_in0[53]),
	.v2c_53_out1 (v2c_in1[53]),
	.v2c_53_out2 (v2c_in2[53]),
	.hard_decision_54 (hard_decision[54]),
	.v2c_54_out0 (v2c_in0[54]),
	.v2c_54_out1 (v2c_in1[54]),
	.v2c_54_out2 (v2c_in2[54]),
	.hard_decision_55 (hard_decision[55]),
	.v2c_55_out0 (v2c_in0[55]),
	.v2c_55_out1 (v2c_in1[55]),
	.v2c_55_out2 (v2c_in2[55]),
	.hard_decision_56 (hard_decision[56]),
	.v2c_56_out0 (v2c_in0[56]),
	.v2c_56_out1 (v2c_in1[56]),
	.v2c_56_out2 (v2c_in2[56]),
	.hard_decision_57 (hard_decision[57]),
	.v2c_57_out0 (v2c_in0[57]),
	.v2c_57_out1 (v2c_in1[57]),
	.v2c_57_out2 (v2c_in2[57]),
	.hard_decision_58 (hard_decision[58]),
	.v2c_58_out0 (v2c_in0[58]),
	.v2c_58_out1 (v2c_in1[58]),
	.v2c_58_out2 (v2c_in2[58]),
	.hard_decision_59 (hard_decision[59]),
	.v2c_59_out0 (v2c_in0[59]),
	.v2c_59_out1 (v2c_in1[59]),
	.v2c_59_out2 (v2c_in2[59]),
	.hard_decision_60 (hard_decision[60]),
	.v2c_60_out0 (v2c_in0[60]),
	.v2c_60_out1 (v2c_in1[60]),
	.v2c_60_out2 (v2c_in2[60]),
	.hard_decision_61 (hard_decision[61]),
	.v2c_61_out0 (v2c_in0[61]),
	.v2c_61_out1 (v2c_in1[61]),
	.v2c_61_out2 (v2c_in2[61]),
	.hard_decision_62 (hard_decision[62]),
	.v2c_62_out0 (v2c_in0[62]),
	.v2c_62_out1 (v2c_in1[62]),
	.v2c_62_out2 (v2c_in2[62]),
	.hard_decision_63 (hard_decision[63]),
	.v2c_63_out0 (v2c_in0[63]),
	.v2c_63_out1 (v2c_in1[63]),
	.v2c_63_out2 (v2c_in2[63]),
	.hard_decision_64 (hard_decision[64]),
	.v2c_64_out0 (v2c_in0[64]),
	.v2c_64_out1 (v2c_in1[64]),
	.v2c_64_out2 (v2c_in2[64]),
	.hard_decision_65 (hard_decision[65]),
	.v2c_65_out0 (v2c_in0[65]),
	.v2c_65_out1 (v2c_in1[65]),
	.v2c_65_out2 (v2c_in2[65]),
	.hard_decision_66 (hard_decision[66]),
	.v2c_66_out0 (v2c_in0[66]),
	.v2c_66_out1 (v2c_in1[66]),
	.v2c_66_out2 (v2c_in2[66]),
	.hard_decision_67 (hard_decision[67]),
	.v2c_67_out0 (v2c_in0[67]),
	.v2c_67_out1 (v2c_in1[67]),
	.v2c_67_out2 (v2c_in2[67]),
	.hard_decision_68 (hard_decision[68]),
	.v2c_68_out0 (v2c_in0[68]),
	.v2c_68_out1 (v2c_in1[68]),
	.v2c_68_out2 (v2c_in2[68]),
	.hard_decision_69 (hard_decision[69]),
	.v2c_69_out0 (v2c_in0[69]),
	.v2c_69_out1 (v2c_in1[69]),
	.v2c_69_out2 (v2c_in2[69]),
	.hard_decision_70 (hard_decision[70]),
	.v2c_70_out0 (v2c_in0[70]),
	.v2c_70_out1 (v2c_in1[70]),
	.v2c_70_out2 (v2c_in2[70]),
	.hard_decision_71 (hard_decision[71]),
	.v2c_71_out0 (v2c_in0[71]),
	.v2c_71_out1 (v2c_in1[71]),
	.v2c_71_out2 (v2c_in2[71]),
	.hard_decision_72 (hard_decision[72]),
	.v2c_72_out0 (v2c_in0[72]),
	.v2c_72_out1 (v2c_in1[72]),
	.v2c_72_out2 (v2c_in2[72]),
	.hard_decision_73 (hard_decision[73]),
	.v2c_73_out0 (v2c_in0[73]),
	.v2c_73_out1 (v2c_in1[73]),
	.v2c_73_out2 (v2c_in2[73]),
	.hard_decision_74 (hard_decision[74]),
	.v2c_74_out0 (v2c_in0[74]),
	.v2c_74_out1 (v2c_in1[74]),
	.v2c_74_out2 (v2c_in2[74]),
	.hard_decision_75 (hard_decision[75]),
	.v2c_75_out0 (v2c_in0[75]),
	.v2c_75_out1 (v2c_in1[75]),
	.v2c_75_out2 (v2c_in2[75]),
	.hard_decision_76 (hard_decision[76]),
	.v2c_76_out0 (v2c_in0[76]),
	.v2c_76_out1 (v2c_in1[76]),
	.v2c_76_out2 (v2c_in2[76]),
	.hard_decision_77 (hard_decision[77]),
	.v2c_77_out0 (v2c_in0[77]),
	.v2c_77_out1 (v2c_in1[77]),
	.v2c_77_out2 (v2c_in2[77]),
	.hard_decision_78 (hard_decision[78]),
	.v2c_78_out0 (v2c_in0[78]),
	.v2c_78_out1 (v2c_in1[78]),
	.v2c_78_out2 (v2c_in2[78]),
	.hard_decision_79 (hard_decision[79]),
	.v2c_79_out0 (v2c_in0[79]),
	.v2c_79_out1 (v2c_in1[79]),
	.v2c_79_out2 (v2c_in2[79]),
	.hard_decision_80 (hard_decision[80]),
	.v2c_80_out0 (v2c_in0[80]),
	.v2c_80_out1 (v2c_in1[80]),
	.v2c_80_out2 (v2c_in2[80]),
	.hard_decision_81 (hard_decision[81]),
	.v2c_81_out0 (v2c_in0[81]),
	.v2c_81_out1 (v2c_in1[81]),
	.v2c_81_out2 (v2c_in2[81]),
	.hard_decision_82 (hard_decision[82]),
	.v2c_82_out0 (v2c_in0[82]),
	.v2c_82_out1 (v2c_in1[82]),
	.v2c_82_out2 (v2c_in2[82]),
	.hard_decision_83 (hard_decision[83]),
	.v2c_83_out0 (v2c_in0[83]),
	.v2c_83_out1 (v2c_in1[83]),
	.v2c_83_out2 (v2c_in2[83]),
	.hard_decision_84 (hard_decision[84]),
	.v2c_84_out0 (v2c_in0[84]),
	.v2c_84_out1 (v2c_in1[84]),
	.v2c_84_out2 (v2c_in2[84]),
	.hard_decision_85 (hard_decision[85]),
	.v2c_85_out0 (v2c_in0[85]),
	.v2c_85_out1 (v2c_in1[85]),
	.v2c_85_out2 (v2c_in2[85]),
	.hard_decision_86 (hard_decision[86]),
	.v2c_86_out0 (v2c_in0[86]),
	.v2c_86_out1 (v2c_in1[86]),
	.v2c_86_out2 (v2c_in2[86]),
	.hard_decision_87 (hard_decision[87]),
	.v2c_87_out0 (v2c_in0[87]),
	.v2c_87_out1 (v2c_in1[87]),
	.v2c_87_out2 (v2c_in2[87]),
	.hard_decision_88 (hard_decision[88]),
	.v2c_88_out0 (v2c_in0[88]),
	.v2c_88_out1 (v2c_in1[88]),
	.v2c_88_out2 (v2c_in2[88]),
	.hard_decision_89 (hard_decision[89]),
	.v2c_89_out0 (v2c_in0[89]),
	.v2c_89_out1 (v2c_in1[89]),
	.v2c_89_out2 (v2c_in2[89]),
	.hard_decision_90 (hard_decision[90]),
	.v2c_90_out0 (v2c_in0[90]),
	.v2c_90_out1 (v2c_in1[90]),
	.v2c_90_out2 (v2c_in2[90]),
	.hard_decision_91 (hard_decision[91]),
	.v2c_91_out0 (v2c_in0[91]),
	.v2c_91_out1 (v2c_in1[91]),
	.v2c_91_out2 (v2c_in2[91]),
	.hard_decision_92 (hard_decision[92]),
	.v2c_92_out0 (v2c_in0[92]),
	.v2c_92_out1 (v2c_in1[92]),
	.v2c_92_out2 (v2c_in2[92]),
	.hard_decision_93 (hard_decision[93]),
	.v2c_93_out0 (v2c_in0[93]),
	.v2c_93_out1 (v2c_in1[93]),
	.v2c_93_out2 (v2c_in2[93]),
	.hard_decision_94 (hard_decision[94]),
	.v2c_94_out0 (v2c_in0[94]),
	.v2c_94_out1 (v2c_in1[94]),
	.v2c_94_out2 (v2c_in2[94]),
	.hard_decision_95 (hard_decision[95]),
	.v2c_95_out0 (v2c_in0[95]),
	.v2c_95_out1 (v2c_in1[95]),
	.v2c_95_out2 (v2c_in2[95]),
	.hard_decision_96 (hard_decision[96]),
	.v2c_96_out0 (v2c_in0[96]),
	.v2c_96_out1 (v2c_in1[96]),
	.v2c_96_out2 (v2c_in2[96]),
	.hard_decision_97 (hard_decision[97]),
	.v2c_97_out0 (v2c_in0[97]),
	.v2c_97_out1 (v2c_in1[97]),
	.v2c_97_out2 (v2c_in2[97]),
	.hard_decision_98 (hard_decision[98]),
	.v2c_98_out0 (v2c_in0[98]),
	.v2c_98_out1 (v2c_in1[98]),
	.v2c_98_out2 (v2c_in2[98]),
	.hard_decision_99 (hard_decision[99]),
	.v2c_99_out0 (v2c_in0[99]),
	.v2c_99_out1 (v2c_in1[99]),
	.v2c_99_out2 (v2c_in2[99]),
	.hard_decision_100 (hard_decision[100]),
	.v2c_100_out0 (v2c_in0[100]),
	.v2c_100_out1 (v2c_in1[100]),
	.v2c_100_out2 (v2c_in2[100]),
	.hard_decision_101 (hard_decision[101]),
	.v2c_101_out0 (v2c_in0[101]),
	.v2c_101_out1 (v2c_in1[101]),
	.v2c_101_out2 (v2c_in2[101]),
	.hard_decision_102 (hard_decision[102]),
	.v2c_102_out0 (v2c_in0[102]),
	.v2c_102_out1 (v2c_in1[102]),
	.v2c_102_out2 (v2c_in2[102]),
	.hard_decision_103 (hard_decision[103]),
	.v2c_103_out0 (v2c_in0[103]),
	.v2c_103_out1 (v2c_in1[103]),
	.v2c_103_out2 (v2c_in2[103]),
	.hard_decision_104 (hard_decision[104]),
	.v2c_104_out0 (v2c_in0[104]),
	.v2c_104_out1 (v2c_in1[104]),
	.v2c_104_out2 (v2c_in2[104]),
	.hard_decision_105 (hard_decision[105]),
	.v2c_105_out0 (v2c_in0[105]),
	.v2c_105_out1 (v2c_in1[105]),
	.v2c_105_out2 (v2c_in2[105]),
	.hard_decision_106 (hard_decision[106]),
	.v2c_106_out0 (v2c_in0[106]),
	.v2c_106_out1 (v2c_in1[106]),
	.v2c_106_out2 (v2c_in2[106]),
	.hard_decision_107 (hard_decision[107]),
	.v2c_107_out0 (v2c_in0[107]),
	.v2c_107_out1 (v2c_in1[107]),
	.v2c_107_out2 (v2c_in2[107]),
	.hard_decision_108 (hard_decision[108]),
	.v2c_108_out0 (v2c_in0[108]),
	.v2c_108_out1 (v2c_in1[108]),
	.v2c_108_out2 (v2c_in2[108]),
	.hard_decision_109 (hard_decision[109]),
	.v2c_109_out0 (v2c_in0[109]),
	.v2c_109_out1 (v2c_in1[109]),
	.v2c_109_out2 (v2c_in2[109]),
	.hard_decision_110 (hard_decision[110]),
	.v2c_110_out0 (v2c_in0[110]),
	.v2c_110_out1 (v2c_in1[110]),
	.v2c_110_out2 (v2c_in2[110]),
	.hard_decision_111 (hard_decision[111]),
	.v2c_111_out0 (v2c_in0[111]),
	.v2c_111_out1 (v2c_in1[111]),
	.v2c_111_out2 (v2c_in2[111]),
	.hard_decision_112 (hard_decision[112]),
	.v2c_112_out0 (v2c_in0[112]),
	.v2c_112_out1 (v2c_in1[112]),
	.v2c_112_out2 (v2c_in2[112]),
	.hard_decision_113 (hard_decision[113]),
	.v2c_113_out0 (v2c_in0[113]),
	.v2c_113_out1 (v2c_in1[113]),
	.v2c_113_out2 (v2c_in2[113]),
	.hard_decision_114 (hard_decision[114]),
	.v2c_114_out0 (v2c_in0[114]),
	.v2c_114_out1 (v2c_in1[114]),
	.v2c_114_out2 (v2c_in2[114]),
	.hard_decision_115 (hard_decision[115]),
	.v2c_115_out0 (v2c_in0[115]),
	.v2c_115_out1 (v2c_in1[115]),
	.v2c_115_out2 (v2c_in2[115]),
	.hard_decision_116 (hard_decision[116]),
	.v2c_116_out0 (v2c_in0[116]),
	.v2c_116_out1 (v2c_in1[116]),
	.v2c_116_out2 (v2c_in2[116]),
	.hard_decision_117 (hard_decision[117]),
	.v2c_117_out0 (v2c_in0[117]),
	.v2c_117_out1 (v2c_in1[117]),
	.v2c_117_out2 (v2c_in2[117]),
	.hard_decision_118 (hard_decision[118]),
	.v2c_118_out0 (v2c_in0[118]),
	.v2c_118_out1 (v2c_in1[118]),
	.v2c_118_out2 (v2c_in2[118]),
	.hard_decision_119 (hard_decision[119]),
	.v2c_119_out0 (v2c_in0[119]),
	.v2c_119_out1 (v2c_in1[119]),
	.v2c_119_out2 (v2c_in2[119]),
	.hard_decision_120 (hard_decision[120]),
	.v2c_120_out0 (v2c_in0[120]),
	.v2c_120_out1 (v2c_in1[120]),
	.v2c_120_out2 (v2c_in2[120]),
	.hard_decision_121 (hard_decision[121]),
	.v2c_121_out0 (v2c_in0[121]),
	.v2c_121_out1 (v2c_in1[121]),
	.v2c_121_out2 (v2c_in2[121]),
	.hard_decision_122 (hard_decision[122]),
	.v2c_122_out0 (v2c_in0[122]),
	.v2c_122_out1 (v2c_in1[122]),
	.v2c_122_out2 (v2c_in2[122]),
	.hard_decision_123 (hard_decision[123]),
	.v2c_123_out0 (v2c_in0[123]),
	.v2c_123_out1 (v2c_in1[123]),
	.v2c_123_out2 (v2c_in2[123]),
	.hard_decision_124 (hard_decision[124]),
	.v2c_124_out0 (v2c_in0[124]),
	.v2c_124_out1 (v2c_in1[124]),
	.v2c_124_out2 (v2c_in2[124]),
	.hard_decision_125 (hard_decision[125]),
	.v2c_125_out0 (v2c_in0[125]),
	.v2c_125_out1 (v2c_in1[125]),
	.v2c_125_out2 (v2c_in2[125]),
	.hard_decision_126 (hard_decision[126]),
	.v2c_126_out0 (v2c_in0[126]),
	.v2c_126_out1 (v2c_in1[126]),
	.v2c_126_out2 (v2c_in2[126]),
	.hard_decision_127 (hard_decision[127]),
	.v2c_127_out0 (v2c_in0[127]),
	.v2c_127_out1 (v2c_in1[127]),
	.v2c_127_out2 (v2c_in2[127]),
	.hard_decision_128 (hard_decision[128]),
	.v2c_128_out0 (v2c_in0[128]),
	.v2c_128_out1 (v2c_in1[128]),
	.v2c_128_out2 (v2c_in2[128]),
	.hard_decision_129 (hard_decision[129]),
	.v2c_129_out0 (v2c_in0[129]),
	.v2c_129_out1 (v2c_in1[129]),
	.v2c_129_out2 (v2c_in2[129]),
	.hard_decision_130 (hard_decision[130]),
	.v2c_130_out0 (v2c_in0[130]),
	.v2c_130_out1 (v2c_in1[130]),
	.v2c_130_out2 (v2c_in2[130]),
	.hard_decision_131 (hard_decision[131]),
	.v2c_131_out0 (v2c_in0[131]),
	.v2c_131_out1 (v2c_in1[131]),
	.v2c_131_out2 (v2c_in2[131]),
	.hard_decision_132 (hard_decision[132]),
	.v2c_132_out0 (v2c_in0[132]),
	.v2c_132_out1 (v2c_in1[132]),
	.v2c_132_out2 (v2c_in2[132]),
	.hard_decision_133 (hard_decision[133]),
	.v2c_133_out0 (v2c_in0[133]),
	.v2c_133_out1 (v2c_in1[133]),
	.v2c_133_out2 (v2c_in2[133]),
	.hard_decision_134 (hard_decision[134]),
	.v2c_134_out0 (v2c_in0[134]),
	.v2c_134_out1 (v2c_in1[134]),
	.v2c_134_out2 (v2c_in2[134]),
	.hard_decision_135 (hard_decision[135]),
	.v2c_135_out0 (v2c_in0[135]),
	.v2c_135_out1 (v2c_in1[135]),
	.v2c_135_out2 (v2c_in2[135]),
	.hard_decision_136 (hard_decision[136]),
	.v2c_136_out0 (v2c_in0[136]),
	.v2c_136_out1 (v2c_in1[136]),
	.v2c_136_out2 (v2c_in2[136]),
	.hard_decision_137 (hard_decision[137]),
	.v2c_137_out0 (v2c_in0[137]),
	.v2c_137_out1 (v2c_in1[137]),
	.v2c_137_out2 (v2c_in2[137]),
	.hard_decision_138 (hard_decision[138]),
	.v2c_138_out0 (v2c_in0[138]),
	.v2c_138_out1 (v2c_in1[138]),
	.v2c_138_out2 (v2c_in2[138]),
	.hard_decision_139 (hard_decision[139]),
	.v2c_139_out0 (v2c_in0[139]),
	.v2c_139_out1 (v2c_in1[139]),
	.v2c_139_out2 (v2c_in2[139]),
	.hard_decision_140 (hard_decision[140]),
	.v2c_140_out0 (v2c_in0[140]),
	.v2c_140_out1 (v2c_in1[140]),
	.v2c_140_out2 (v2c_in2[140]),
	.hard_decision_141 (hard_decision[141]),
	.v2c_141_out0 (v2c_in0[141]),
	.v2c_141_out1 (v2c_in1[141]),
	.v2c_141_out2 (v2c_in2[141]),
	.hard_decision_142 (hard_decision[142]),
	.v2c_142_out0 (v2c_in0[142]),
	.v2c_142_out1 (v2c_in1[142]),
	.v2c_142_out2 (v2c_in2[142]),
	.hard_decision_143 (hard_decision[143]),
	.v2c_143_out0 (v2c_in0[143]),
	.v2c_143_out1 (v2c_in1[143]),
	.v2c_143_out2 (v2c_in2[143]),
	.hard_decision_144 (hard_decision[144]),
	.v2c_144_out0 (v2c_in0[144]),
	.v2c_144_out1 (v2c_in1[144]),
	.v2c_144_out2 (v2c_in2[144]),
	.hard_decision_145 (hard_decision[145]),
	.v2c_145_out0 (v2c_in0[145]),
	.v2c_145_out1 (v2c_in1[145]),
	.v2c_145_out2 (v2c_in2[145]),
	.hard_decision_146 (hard_decision[146]),
	.v2c_146_out0 (v2c_in0[146]),
	.v2c_146_out1 (v2c_in1[146]),
	.v2c_146_out2 (v2c_in2[146]),
	.hard_decision_147 (hard_decision[147]),
	.v2c_147_out0 (v2c_in0[147]),
	.v2c_147_out1 (v2c_in1[147]),
	.v2c_147_out2 (v2c_in2[147]),
	.hard_decision_148 (hard_decision[148]),
	.v2c_148_out0 (v2c_in0[148]),
	.v2c_148_out1 (v2c_in1[148]),
	.v2c_148_out2 (v2c_in2[148]),
	.hard_decision_149 (hard_decision[149]),
	.v2c_149_out0 (v2c_in0[149]),
	.v2c_149_out1 (v2c_in1[149]),
	.v2c_149_out2 (v2c_in2[149]),
	.hard_decision_150 (hard_decision[150]),
	.v2c_150_out0 (v2c_in0[150]),
	.v2c_150_out1 (v2c_in1[150]),
	.v2c_150_out2 (v2c_in2[150]),
	.hard_decision_151 (hard_decision[151]),
	.v2c_151_out0 (v2c_in0[151]),
	.v2c_151_out1 (v2c_in1[151]),
	.v2c_151_out2 (v2c_in2[151]),
	.hard_decision_152 (hard_decision[152]),
	.v2c_152_out0 (v2c_in0[152]),
	.v2c_152_out1 (v2c_in1[152]),
	.v2c_152_out2 (v2c_in2[152]),
	.hard_decision_153 (hard_decision[153]),
	.v2c_153_out0 (v2c_in0[153]),
	.v2c_153_out1 (v2c_in1[153]),
	.v2c_153_out2 (v2c_in2[153]),
	.hard_decision_154 (hard_decision[154]),
	.v2c_154_out0 (v2c_in0[154]),
	.v2c_154_out1 (v2c_in1[154]),
	.v2c_154_out2 (v2c_in2[154]),
	.hard_decision_155 (hard_decision[155]),
	.v2c_155_out0 (v2c_in0[155]),
	.v2c_155_out1 (v2c_in1[155]),
	.v2c_155_out2 (v2c_in2[155]),
	.hard_decision_156 (hard_decision[156]),
	.v2c_156_out0 (v2c_in0[156]),
	.v2c_156_out1 (v2c_in1[156]),
	.v2c_156_out2 (v2c_in2[156]),
	.hard_decision_157 (hard_decision[157]),
	.v2c_157_out0 (v2c_in0[157]),
	.v2c_157_out1 (v2c_in1[157]),
	.v2c_157_out2 (v2c_in2[157]),
	.hard_decision_158 (hard_decision[158]),
	.v2c_158_out0 (v2c_in0[158]),
	.v2c_158_out1 (v2c_in1[158]),
	.v2c_158_out2 (v2c_in2[158]),
	.hard_decision_159 (hard_decision[159]),
	.v2c_159_out0 (v2c_in0[159]),
	.v2c_159_out1 (v2c_in1[159]),
	.v2c_159_out2 (v2c_in2[159]),
	.hard_decision_160 (hard_decision[160]),
	.v2c_160_out0 (v2c_in0[160]),
	.v2c_160_out1 (v2c_in1[160]),
	.v2c_160_out2 (v2c_in2[160]),
	.hard_decision_161 (hard_decision[161]),
	.v2c_161_out0 (v2c_in0[161]),
	.v2c_161_out1 (v2c_in1[161]),
	.v2c_161_out2 (v2c_in2[161]),
	.hard_decision_162 (hard_decision[162]),
	.v2c_162_out0 (v2c_in0[162]),
	.v2c_162_out1 (v2c_in1[162]),
	.v2c_162_out2 (v2c_in2[162]),
	.hard_decision_163 (hard_decision[163]),
	.v2c_163_out0 (v2c_in0[163]),
	.v2c_163_out1 (v2c_in1[163]),
	.v2c_163_out2 (v2c_in2[163]),
	.hard_decision_164 (hard_decision[164]),
	.v2c_164_out0 (v2c_in0[164]),
	.v2c_164_out1 (v2c_in1[164]),
	.v2c_164_out2 (v2c_in2[164]),
	.hard_decision_165 (hard_decision[165]),
	.v2c_165_out0 (v2c_in0[165]),
	.v2c_165_out1 (v2c_in1[165]),
	.v2c_165_out2 (v2c_in2[165]),
	.hard_decision_166 (hard_decision[166]),
	.v2c_166_out0 (v2c_in0[166]),
	.v2c_166_out1 (v2c_in1[166]),
	.v2c_166_out2 (v2c_in2[166]),
	.hard_decision_167 (hard_decision[167]),
	.v2c_167_out0 (v2c_in0[167]),
	.v2c_167_out1 (v2c_in1[167]),
	.v2c_167_out2 (v2c_in2[167]),
	.hard_decision_168 (hard_decision[168]),
	.v2c_168_out0 (v2c_in0[168]),
	.v2c_168_out1 (v2c_in1[168]),
	.v2c_168_out2 (v2c_in2[168]),
	.hard_decision_169 (hard_decision[169]),
	.v2c_169_out0 (v2c_in0[169]),
	.v2c_169_out1 (v2c_in1[169]),
	.v2c_169_out2 (v2c_in2[169]),
	.hard_decision_170 (hard_decision[170]),
	.v2c_170_out0 (v2c_in0[170]),
	.v2c_170_out1 (v2c_in1[170]),
	.v2c_170_out2 (v2c_in2[170]),
	.hard_decision_171 (hard_decision[171]),
	.v2c_171_out0 (v2c_in0[171]),
	.v2c_171_out1 (v2c_in1[171]),
	.v2c_171_out2 (v2c_in2[171]),
	.hard_decision_172 (hard_decision[172]),
	.v2c_172_out0 (v2c_in0[172]),
	.v2c_172_out1 (v2c_in1[172]),
	.v2c_172_out2 (v2c_in2[172]),
	.hard_decision_173 (hard_decision[173]),
	.v2c_173_out0 (v2c_in0[173]),
	.v2c_173_out1 (v2c_in1[173]),
	.v2c_173_out2 (v2c_in2[173]),
	.hard_decision_174 (hard_decision[174]),
	.v2c_174_out0 (v2c_in0[174]),
	.v2c_174_out1 (v2c_in1[174]),
	.v2c_174_out2 (v2c_in2[174]),
	.hard_decision_175 (hard_decision[175]),
	.v2c_175_out0 (v2c_in0[175]),
	.v2c_175_out1 (v2c_in1[175]),
	.v2c_175_out2 (v2c_in2[175]),
	.hard_decision_176 (hard_decision[176]),
	.v2c_176_out0 (v2c_in0[176]),
	.v2c_176_out1 (v2c_in1[176]),
	.v2c_176_out2 (v2c_in2[176]),
	.hard_decision_177 (hard_decision[177]),
	.v2c_177_out0 (v2c_in0[177]),
	.v2c_177_out1 (v2c_in1[177]),
	.v2c_177_out2 (v2c_in2[177]),
	.hard_decision_178 (hard_decision[178]),
	.v2c_178_out0 (v2c_in0[178]),
	.v2c_178_out1 (v2c_in1[178]),
	.v2c_178_out2 (v2c_in2[178]),
	.hard_decision_179 (hard_decision[179]),
	.v2c_179_out0 (v2c_in0[179]),
	.v2c_179_out1 (v2c_in1[179]),
	.v2c_179_out2 (v2c_in2[179]),
	.hard_decision_180 (hard_decision[180]),
	.v2c_180_out0 (v2c_in0[180]),
	.v2c_180_out1 (v2c_in1[180]),
	.v2c_180_out2 (v2c_in2[180]),
	.hard_decision_181 (hard_decision[181]),
	.v2c_181_out0 (v2c_in0[181]),
	.v2c_181_out1 (v2c_in1[181]),
	.v2c_181_out2 (v2c_in2[181]),
	.hard_decision_182 (hard_decision[182]),
	.v2c_182_out0 (v2c_in0[182]),
	.v2c_182_out1 (v2c_in1[182]),
	.v2c_182_out2 (v2c_in2[182]),
	.hard_decision_183 (hard_decision[183]),
	.v2c_183_out0 (v2c_in0[183]),
	.v2c_183_out1 (v2c_in1[183]),
	.v2c_183_out2 (v2c_in2[183]),
	.hard_decision_184 (hard_decision[184]),
	.v2c_184_out0 (v2c_in0[184]),
	.v2c_184_out1 (v2c_in1[184]),
	.v2c_184_out2 (v2c_in2[184]),
	.hard_decision_185 (hard_decision[185]),
	.v2c_185_out0 (v2c_in0[185]),
	.v2c_185_out1 (v2c_in1[185]),
	.v2c_185_out2 (v2c_in2[185]),
	.hard_decision_186 (hard_decision[186]),
	.v2c_186_out0 (v2c_in0[186]),
	.v2c_186_out1 (v2c_in1[186]),
	.v2c_186_out2 (v2c_in2[186]),
	.hard_decision_187 (hard_decision[187]),
	.v2c_187_out0 (v2c_in0[187]),
	.v2c_187_out1 (v2c_in1[187]),
	.v2c_187_out2 (v2c_in2[187]),
	.hard_decision_188 (hard_decision[188]),
	.v2c_188_out0 (v2c_in0[188]),
	.v2c_188_out1 (v2c_in1[188]),
	.v2c_188_out2 (v2c_in2[188]),
	.hard_decision_189 (hard_decision[189]),
	.v2c_189_out0 (v2c_in0[189]),
	.v2c_189_out1 (v2c_in1[189]),
	.v2c_189_out2 (v2c_in2[189]),
	.hard_decision_190 (hard_decision[190]),
	.v2c_190_out0 (v2c_in0[190]),
	.v2c_190_out1 (v2c_in1[190]),
	.v2c_190_out2 (v2c_in2[190]),
	.hard_decision_191 (hard_decision[191]),
	.v2c_191_out0 (v2c_in0[191]),
	.v2c_191_out1 (v2c_in1[191]),
	.v2c_191_out2 (v2c_in2[191]),
	.hard_decision_192 (hard_decision[192]),
	.v2c_192_out0 (v2c_in0[192]),
	.v2c_192_out1 (v2c_in1[192]),
	.v2c_192_out2 (v2c_in2[192]),
	.hard_decision_193 (hard_decision[193]),
	.v2c_193_out0 (v2c_in0[193]),
	.v2c_193_out1 (v2c_in1[193]),
	.v2c_193_out2 (v2c_in2[193]),
	.hard_decision_194 (hard_decision[194]),
	.v2c_194_out0 (v2c_in0[194]),
	.v2c_194_out1 (v2c_in1[194]),
	.v2c_194_out2 (v2c_in2[194]),
	.hard_decision_195 (hard_decision[195]),
	.v2c_195_out0 (v2c_in0[195]),
	.v2c_195_out1 (v2c_in1[195]),
	.v2c_195_out2 (v2c_in2[195]),
	.hard_decision_196 (hard_decision[196]),
	.v2c_196_out0 (v2c_in0[196]),
	.v2c_196_out1 (v2c_in1[196]),
	.v2c_196_out2 (v2c_in2[196]),
	.hard_decision_197 (hard_decision[197]),
	.v2c_197_out0 (v2c_in0[197]),
	.v2c_197_out1 (v2c_in1[197]),
	.v2c_197_out2 (v2c_in2[197]),
	.hard_decision_198 (hard_decision[198]),
	.v2c_198_out0 (v2c_in0[198]),
	.v2c_198_out1 (v2c_in1[198]),
	.v2c_198_out2 (v2c_in2[198]),
	.hard_decision_199 (hard_decision[199]),
	.v2c_199_out0 (v2c_in0[199]),
	.v2c_199_out1 (v2c_in1[199]),
	.v2c_199_out2 (v2c_in2[199]),
	.hard_decision_200 (hard_decision[200]),
	.v2c_200_out0 (v2c_in0[200]),
	.v2c_200_out1 (v2c_in1[200]),
	.v2c_200_out2 (v2c_in2[200]),
	.hard_decision_201 (hard_decision[201]),
	.v2c_201_out0 (v2c_in0[201]),
	.v2c_201_out1 (v2c_in1[201]),
	.v2c_201_out2 (v2c_in2[201]),
	.hard_decision_202 (hard_decision[202]),
	.v2c_202_out0 (v2c_in0[202]),
	.v2c_202_out1 (v2c_in1[202]),
	.v2c_202_out2 (v2c_in2[202]),
	.hard_decision_203 (hard_decision[203]),
	.v2c_203_out0 (v2c_in0[203]),
	.v2c_203_out1 (v2c_in1[203]),
	.v2c_203_out2 (v2c_in2[203]),

	.ch_msg_0 (ch_msg_0[DATAPATH_WIDTH-1:0]),
	.c2v_0_in0 (c2v_out0[0]),
	.c2v_0_in1 (c2v_out1[0]),
	.c2v_0_in2 (c2v_out2[0]),
	.ch_msg_1 (ch_msg_1[DATAPATH_WIDTH-1:0]),
	.c2v_1_in0 (c2v_out0[1]),
	.c2v_1_in1 (c2v_out1[1]),
	.c2v_1_in2 (c2v_out2[1]),
	.ch_msg_2 (ch_msg_2[DATAPATH_WIDTH-1:0]),
	.c2v_2_in0 (c2v_out0[2]),
	.c2v_2_in1 (c2v_out1[2]),
	.c2v_2_in2 (c2v_out2[2]),
	.ch_msg_3 (ch_msg_3[DATAPATH_WIDTH-1:0]),
	.c2v_3_in0 (c2v_out0[3]),
	.c2v_3_in1 (c2v_out1[3]),
	.c2v_3_in2 (c2v_out2[3]),
	.ch_msg_4 (ch_msg_4[DATAPATH_WIDTH-1:0]),
	.c2v_4_in0 (c2v_out0[4]),
	.c2v_4_in1 (c2v_out1[4]),
	.c2v_4_in2 (c2v_out2[4]),
	.ch_msg_5 (ch_msg_5[DATAPATH_WIDTH-1:0]),
	.c2v_5_in0 (c2v_out0[5]),
	.c2v_5_in1 (c2v_out1[5]),
	.c2v_5_in2 (c2v_out2[5]),
	.ch_msg_6 (ch_msg_6[DATAPATH_WIDTH-1:0]),
	.c2v_6_in0 (c2v_out0[6]),
	.c2v_6_in1 (c2v_out1[6]),
	.c2v_6_in2 (c2v_out2[6]),
	.ch_msg_7 (ch_msg_7[DATAPATH_WIDTH-1:0]),
	.c2v_7_in0 (c2v_out0[7]),
	.c2v_7_in1 (c2v_out1[7]),
	.c2v_7_in2 (c2v_out2[7]),
	.ch_msg_8 (ch_msg_8[DATAPATH_WIDTH-1:0]),
	.c2v_8_in0 (c2v_out0[8]),
	.c2v_8_in1 (c2v_out1[8]),
	.c2v_8_in2 (c2v_out2[8]),
	.ch_msg_9 (ch_msg_9[DATAPATH_WIDTH-1:0]),
	.c2v_9_in0 (c2v_out0[9]),
	.c2v_9_in1 (c2v_out1[9]),
	.c2v_9_in2 (c2v_out2[9]),
	.ch_msg_10 (ch_msg_10[DATAPATH_WIDTH-1:0]),
	.c2v_10_in0 (c2v_out0[10]),
	.c2v_10_in1 (c2v_out1[10]),
	.c2v_10_in2 (c2v_out2[10]),
	.ch_msg_11 (ch_msg_11[DATAPATH_WIDTH-1:0]),
	.c2v_11_in0 (c2v_out0[11]),
	.c2v_11_in1 (c2v_out1[11]),
	.c2v_11_in2 (c2v_out2[11]),
	.ch_msg_12 (ch_msg_12[DATAPATH_WIDTH-1:0]),
	.c2v_12_in0 (c2v_out0[12]),
	.c2v_12_in1 (c2v_out1[12]),
	.c2v_12_in2 (c2v_out2[12]),
	.ch_msg_13 (ch_msg_13[DATAPATH_WIDTH-1:0]),
	.c2v_13_in0 (c2v_out0[13]),
	.c2v_13_in1 (c2v_out1[13]),
	.c2v_13_in2 (c2v_out2[13]),
	.ch_msg_14 (ch_msg_14[DATAPATH_WIDTH-1:0]),
	.c2v_14_in0 (c2v_out0[14]),
	.c2v_14_in1 (c2v_out1[14]),
	.c2v_14_in2 (c2v_out2[14]),
	.ch_msg_15 (ch_msg_15[DATAPATH_WIDTH-1:0]),
	.c2v_15_in0 (c2v_out0[15]),
	.c2v_15_in1 (c2v_out1[15]),
	.c2v_15_in2 (c2v_out2[15]),
	.ch_msg_16 (ch_msg_16[DATAPATH_WIDTH-1:0]),
	.c2v_16_in0 (c2v_out0[16]),
	.c2v_16_in1 (c2v_out1[16]),
	.c2v_16_in2 (c2v_out2[16]),
	.ch_msg_17 (ch_msg_17[DATAPATH_WIDTH-1:0]),
	.c2v_17_in0 (c2v_out0[17]),
	.c2v_17_in1 (c2v_out1[17]),
	.c2v_17_in2 (c2v_out2[17]),
	.ch_msg_18 (ch_msg_18[DATAPATH_WIDTH-1:0]),
	.c2v_18_in0 (c2v_out0[18]),
	.c2v_18_in1 (c2v_out1[18]),
	.c2v_18_in2 (c2v_out2[18]),
	.ch_msg_19 (ch_msg_19[DATAPATH_WIDTH-1:0]),
	.c2v_19_in0 (c2v_out0[19]),
	.c2v_19_in1 (c2v_out1[19]),
	.c2v_19_in2 (c2v_out2[19]),
	.ch_msg_20 (ch_msg_20[DATAPATH_WIDTH-1:0]),
	.c2v_20_in0 (c2v_out0[20]),
	.c2v_20_in1 (c2v_out1[20]),
	.c2v_20_in2 (c2v_out2[20]),
	.ch_msg_21 (ch_msg_21[DATAPATH_WIDTH-1:0]),
	.c2v_21_in0 (c2v_out0[21]),
	.c2v_21_in1 (c2v_out1[21]),
	.c2v_21_in2 (c2v_out2[21]),
	.ch_msg_22 (ch_msg_22[DATAPATH_WIDTH-1:0]),
	.c2v_22_in0 (c2v_out0[22]),
	.c2v_22_in1 (c2v_out1[22]),
	.c2v_22_in2 (c2v_out2[22]),
	.ch_msg_23 (ch_msg_23[DATAPATH_WIDTH-1:0]),
	.c2v_23_in0 (c2v_out0[23]),
	.c2v_23_in1 (c2v_out1[23]),
	.c2v_23_in2 (c2v_out2[23]),
	.ch_msg_24 (ch_msg_24[DATAPATH_WIDTH-1:0]),
	.c2v_24_in0 (c2v_out0[24]),
	.c2v_24_in1 (c2v_out1[24]),
	.c2v_24_in2 (c2v_out2[24]),
	.ch_msg_25 (ch_msg_25[DATAPATH_WIDTH-1:0]),
	.c2v_25_in0 (c2v_out0[25]),
	.c2v_25_in1 (c2v_out1[25]),
	.c2v_25_in2 (c2v_out2[25]),
	.ch_msg_26 (ch_msg_26[DATAPATH_WIDTH-1:0]),
	.c2v_26_in0 (c2v_out0[26]),
	.c2v_26_in1 (c2v_out1[26]),
	.c2v_26_in2 (c2v_out2[26]),
	.ch_msg_27 (ch_msg_27[DATAPATH_WIDTH-1:0]),
	.c2v_27_in0 (c2v_out0[27]),
	.c2v_27_in1 (c2v_out1[27]),
	.c2v_27_in2 (c2v_out2[27]),
	.ch_msg_28 (ch_msg_28[DATAPATH_WIDTH-1:0]),
	.c2v_28_in0 (c2v_out0[28]),
	.c2v_28_in1 (c2v_out1[28]),
	.c2v_28_in2 (c2v_out2[28]),
	.ch_msg_29 (ch_msg_29[DATAPATH_WIDTH-1:0]),
	.c2v_29_in0 (c2v_out0[29]),
	.c2v_29_in1 (c2v_out1[29]),
	.c2v_29_in2 (c2v_out2[29]),
	.ch_msg_30 (ch_msg_30[DATAPATH_WIDTH-1:0]),
	.c2v_30_in0 (c2v_out0[30]),
	.c2v_30_in1 (c2v_out1[30]),
	.c2v_30_in2 (c2v_out2[30]),
	.ch_msg_31 (ch_msg_31[DATAPATH_WIDTH-1:0]),
	.c2v_31_in0 (c2v_out0[31]),
	.c2v_31_in1 (c2v_out1[31]),
	.c2v_31_in2 (c2v_out2[31]),
	.ch_msg_32 (ch_msg_32[DATAPATH_WIDTH-1:0]),
	.c2v_32_in0 (c2v_out0[32]),
	.c2v_32_in1 (c2v_out1[32]),
	.c2v_32_in2 (c2v_out2[32]),
	.ch_msg_33 (ch_msg_33[DATAPATH_WIDTH-1:0]),
	.c2v_33_in0 (c2v_out0[33]),
	.c2v_33_in1 (c2v_out1[33]),
	.c2v_33_in2 (c2v_out2[33]),
	.ch_msg_34 (ch_msg_34[DATAPATH_WIDTH-1:0]),
	.c2v_34_in0 (c2v_out0[34]),
	.c2v_34_in1 (c2v_out1[34]),
	.c2v_34_in2 (c2v_out2[34]),
	.ch_msg_35 (ch_msg_35[DATAPATH_WIDTH-1:0]),
	.c2v_35_in0 (c2v_out0[35]),
	.c2v_35_in1 (c2v_out1[35]),
	.c2v_35_in2 (c2v_out2[35]),
	.ch_msg_36 (ch_msg_36[DATAPATH_WIDTH-1:0]),
	.c2v_36_in0 (c2v_out0[36]),
	.c2v_36_in1 (c2v_out1[36]),
	.c2v_36_in2 (c2v_out2[36]),
	.ch_msg_37 (ch_msg_37[DATAPATH_WIDTH-1:0]),
	.c2v_37_in0 (c2v_out0[37]),
	.c2v_37_in1 (c2v_out1[37]),
	.c2v_37_in2 (c2v_out2[37]),
	.ch_msg_38 (ch_msg_38[DATAPATH_WIDTH-1:0]),
	.c2v_38_in0 (c2v_out0[38]),
	.c2v_38_in1 (c2v_out1[38]),
	.c2v_38_in2 (c2v_out2[38]),
	.ch_msg_39 (ch_msg_39[DATAPATH_WIDTH-1:0]),
	.c2v_39_in0 (c2v_out0[39]),
	.c2v_39_in1 (c2v_out1[39]),
	.c2v_39_in2 (c2v_out2[39]),
	.ch_msg_40 (ch_msg_40[DATAPATH_WIDTH-1:0]),
	.c2v_40_in0 (c2v_out0[40]),
	.c2v_40_in1 (c2v_out1[40]),
	.c2v_40_in2 (c2v_out2[40]),
	.ch_msg_41 (ch_msg_41[DATAPATH_WIDTH-1:0]),
	.c2v_41_in0 (c2v_out0[41]),
	.c2v_41_in1 (c2v_out1[41]),
	.c2v_41_in2 (c2v_out2[41]),
	.ch_msg_42 (ch_msg_42[DATAPATH_WIDTH-1:0]),
	.c2v_42_in0 (c2v_out0[42]),
	.c2v_42_in1 (c2v_out1[42]),
	.c2v_42_in2 (c2v_out2[42]),
	.ch_msg_43 (ch_msg_43[DATAPATH_WIDTH-1:0]),
	.c2v_43_in0 (c2v_out0[43]),
	.c2v_43_in1 (c2v_out1[43]),
	.c2v_43_in2 (c2v_out2[43]),
	.ch_msg_44 (ch_msg_44[DATAPATH_WIDTH-1:0]),
	.c2v_44_in0 (c2v_out0[44]),
	.c2v_44_in1 (c2v_out1[44]),
	.c2v_44_in2 (c2v_out2[44]),
	.ch_msg_45 (ch_msg_45[DATAPATH_WIDTH-1:0]),
	.c2v_45_in0 (c2v_out0[45]),
	.c2v_45_in1 (c2v_out1[45]),
	.c2v_45_in2 (c2v_out2[45]),
	.ch_msg_46 (ch_msg_46[DATAPATH_WIDTH-1:0]),
	.c2v_46_in0 (c2v_out0[46]),
	.c2v_46_in1 (c2v_out1[46]),
	.c2v_46_in2 (c2v_out2[46]),
	.ch_msg_47 (ch_msg_47[DATAPATH_WIDTH-1:0]),
	.c2v_47_in0 (c2v_out0[47]),
	.c2v_47_in1 (c2v_out1[47]),
	.c2v_47_in2 (c2v_out2[47]),
	.ch_msg_48 (ch_msg_48[DATAPATH_WIDTH-1:0]),
	.c2v_48_in0 (c2v_out0[48]),
	.c2v_48_in1 (c2v_out1[48]),
	.c2v_48_in2 (c2v_out2[48]),
	.ch_msg_49 (ch_msg_49[DATAPATH_WIDTH-1:0]),
	.c2v_49_in0 (c2v_out0[49]),
	.c2v_49_in1 (c2v_out1[49]),
	.c2v_49_in2 (c2v_out2[49]),
	.ch_msg_50 (ch_msg_50[DATAPATH_WIDTH-1:0]),
	.c2v_50_in0 (c2v_out0[50]),
	.c2v_50_in1 (c2v_out1[50]),
	.c2v_50_in2 (c2v_out2[50]),
	.ch_msg_51 (ch_msg_51[DATAPATH_WIDTH-1:0]),
	.c2v_51_in0 (c2v_out0[51]),
	.c2v_51_in1 (c2v_out1[51]),
	.c2v_51_in2 (c2v_out2[51]),
	.ch_msg_52 (ch_msg_52[DATAPATH_WIDTH-1:0]),
	.c2v_52_in0 (c2v_out0[52]),
	.c2v_52_in1 (c2v_out1[52]),
	.c2v_52_in2 (c2v_out2[52]),
	.ch_msg_53 (ch_msg_53[DATAPATH_WIDTH-1:0]),
	.c2v_53_in0 (c2v_out0[53]),
	.c2v_53_in1 (c2v_out1[53]),
	.c2v_53_in2 (c2v_out2[53]),
	.ch_msg_54 (ch_msg_54[DATAPATH_WIDTH-1:0]),
	.c2v_54_in0 (c2v_out0[54]),
	.c2v_54_in1 (c2v_out1[54]),
	.c2v_54_in2 (c2v_out2[54]),
	.ch_msg_55 (ch_msg_55[DATAPATH_WIDTH-1:0]),
	.c2v_55_in0 (c2v_out0[55]),
	.c2v_55_in1 (c2v_out1[55]),
	.c2v_55_in2 (c2v_out2[55]),
	.ch_msg_56 (ch_msg_56[DATAPATH_WIDTH-1:0]),
	.c2v_56_in0 (c2v_out0[56]),
	.c2v_56_in1 (c2v_out1[56]),
	.c2v_56_in2 (c2v_out2[56]),
	.ch_msg_57 (ch_msg_57[DATAPATH_WIDTH-1:0]),
	.c2v_57_in0 (c2v_out0[57]),
	.c2v_57_in1 (c2v_out1[57]),
	.c2v_57_in2 (c2v_out2[57]),
	.ch_msg_58 (ch_msg_58[DATAPATH_WIDTH-1:0]),
	.c2v_58_in0 (c2v_out0[58]),
	.c2v_58_in1 (c2v_out1[58]),
	.c2v_58_in2 (c2v_out2[58]),
	.ch_msg_59 (ch_msg_59[DATAPATH_WIDTH-1:0]),
	.c2v_59_in0 (c2v_out0[59]),
	.c2v_59_in1 (c2v_out1[59]),
	.c2v_59_in2 (c2v_out2[59]),
	.ch_msg_60 (ch_msg_60[DATAPATH_WIDTH-1:0]),
	.c2v_60_in0 (c2v_out0[60]),
	.c2v_60_in1 (c2v_out1[60]),
	.c2v_60_in2 (c2v_out2[60]),
	.ch_msg_61 (ch_msg_61[DATAPATH_WIDTH-1:0]),
	.c2v_61_in0 (c2v_out0[61]),
	.c2v_61_in1 (c2v_out1[61]),
	.c2v_61_in2 (c2v_out2[61]),
	.ch_msg_62 (ch_msg_62[DATAPATH_WIDTH-1:0]),
	.c2v_62_in0 (c2v_out0[62]),
	.c2v_62_in1 (c2v_out1[62]),
	.c2v_62_in2 (c2v_out2[62]),
	.ch_msg_63 (ch_msg_63[DATAPATH_WIDTH-1:0]),
	.c2v_63_in0 (c2v_out0[63]),
	.c2v_63_in1 (c2v_out1[63]),
	.c2v_63_in2 (c2v_out2[63]),
	.ch_msg_64 (ch_msg_64[DATAPATH_WIDTH-1:0]),
	.c2v_64_in0 (c2v_out0[64]),
	.c2v_64_in1 (c2v_out1[64]),
	.c2v_64_in2 (c2v_out2[64]),
	.ch_msg_65 (ch_msg_65[DATAPATH_WIDTH-1:0]),
	.c2v_65_in0 (c2v_out0[65]),
	.c2v_65_in1 (c2v_out1[65]),
	.c2v_65_in2 (c2v_out2[65]),
	.ch_msg_66 (ch_msg_66[DATAPATH_WIDTH-1:0]),
	.c2v_66_in0 (c2v_out0[66]),
	.c2v_66_in1 (c2v_out1[66]),
	.c2v_66_in2 (c2v_out2[66]),
	.ch_msg_67 (ch_msg_67[DATAPATH_WIDTH-1:0]),
	.c2v_67_in0 (c2v_out0[67]),
	.c2v_67_in1 (c2v_out1[67]),
	.c2v_67_in2 (c2v_out2[67]),
	.ch_msg_68 (ch_msg_68[DATAPATH_WIDTH-1:0]),
	.c2v_68_in0 (c2v_out0[68]),
	.c2v_68_in1 (c2v_out1[68]),
	.c2v_68_in2 (c2v_out2[68]),
	.ch_msg_69 (ch_msg_69[DATAPATH_WIDTH-1:0]),
	.c2v_69_in0 (c2v_out0[69]),
	.c2v_69_in1 (c2v_out1[69]),
	.c2v_69_in2 (c2v_out2[69]),
	.ch_msg_70 (ch_msg_70[DATAPATH_WIDTH-1:0]),
	.c2v_70_in0 (c2v_out0[70]),
	.c2v_70_in1 (c2v_out1[70]),
	.c2v_70_in2 (c2v_out2[70]),
	.ch_msg_71 (ch_msg_71[DATAPATH_WIDTH-1:0]),
	.c2v_71_in0 (c2v_out0[71]),
	.c2v_71_in1 (c2v_out1[71]),
	.c2v_71_in2 (c2v_out2[71]),
	.ch_msg_72 (ch_msg_72[DATAPATH_WIDTH-1:0]),
	.c2v_72_in0 (c2v_out0[72]),
	.c2v_72_in1 (c2v_out1[72]),
	.c2v_72_in2 (c2v_out2[72]),
	.ch_msg_73 (ch_msg_73[DATAPATH_WIDTH-1:0]),
	.c2v_73_in0 (c2v_out0[73]),
	.c2v_73_in1 (c2v_out1[73]),
	.c2v_73_in2 (c2v_out2[73]),
	.ch_msg_74 (ch_msg_74[DATAPATH_WIDTH-1:0]),
	.c2v_74_in0 (c2v_out0[74]),
	.c2v_74_in1 (c2v_out1[74]),
	.c2v_74_in2 (c2v_out2[74]),
	.ch_msg_75 (ch_msg_75[DATAPATH_WIDTH-1:0]),
	.c2v_75_in0 (c2v_out0[75]),
	.c2v_75_in1 (c2v_out1[75]),
	.c2v_75_in2 (c2v_out2[75]),
	.ch_msg_76 (ch_msg_76[DATAPATH_WIDTH-1:0]),
	.c2v_76_in0 (c2v_out0[76]),
	.c2v_76_in1 (c2v_out1[76]),
	.c2v_76_in2 (c2v_out2[76]),
	.ch_msg_77 (ch_msg_77[DATAPATH_WIDTH-1:0]),
	.c2v_77_in0 (c2v_out0[77]),
	.c2v_77_in1 (c2v_out1[77]),
	.c2v_77_in2 (c2v_out2[77]),
	.ch_msg_78 (ch_msg_78[DATAPATH_WIDTH-1:0]),
	.c2v_78_in0 (c2v_out0[78]),
	.c2v_78_in1 (c2v_out1[78]),
	.c2v_78_in2 (c2v_out2[78]),
	.ch_msg_79 (ch_msg_79[DATAPATH_WIDTH-1:0]),
	.c2v_79_in0 (c2v_out0[79]),
	.c2v_79_in1 (c2v_out1[79]),
	.c2v_79_in2 (c2v_out2[79]),
	.ch_msg_80 (ch_msg_80[DATAPATH_WIDTH-1:0]),
	.c2v_80_in0 (c2v_out0[80]),
	.c2v_80_in1 (c2v_out1[80]),
	.c2v_80_in2 (c2v_out2[80]),
	.ch_msg_81 (ch_msg_81[DATAPATH_WIDTH-1:0]),
	.c2v_81_in0 (c2v_out0[81]),
	.c2v_81_in1 (c2v_out1[81]),
	.c2v_81_in2 (c2v_out2[81]),
	.ch_msg_82 (ch_msg_82[DATAPATH_WIDTH-1:0]),
	.c2v_82_in0 (c2v_out0[82]),
	.c2v_82_in1 (c2v_out1[82]),
	.c2v_82_in2 (c2v_out2[82]),
	.ch_msg_83 (ch_msg_83[DATAPATH_WIDTH-1:0]),
	.c2v_83_in0 (c2v_out0[83]),
	.c2v_83_in1 (c2v_out1[83]),
	.c2v_83_in2 (c2v_out2[83]),
	.ch_msg_84 (ch_msg_84[DATAPATH_WIDTH-1:0]),
	.c2v_84_in0 (c2v_out0[84]),
	.c2v_84_in1 (c2v_out1[84]),
	.c2v_84_in2 (c2v_out2[84]),
	.ch_msg_85 (ch_msg_85[DATAPATH_WIDTH-1:0]),
	.c2v_85_in0 (c2v_out0[85]),
	.c2v_85_in1 (c2v_out1[85]),
	.c2v_85_in2 (c2v_out2[85]),
	.ch_msg_86 (ch_msg_86[DATAPATH_WIDTH-1:0]),
	.c2v_86_in0 (c2v_out0[86]),
	.c2v_86_in1 (c2v_out1[86]),
	.c2v_86_in2 (c2v_out2[86]),
	.ch_msg_87 (ch_msg_87[DATAPATH_WIDTH-1:0]),
	.c2v_87_in0 (c2v_out0[87]),
	.c2v_87_in1 (c2v_out1[87]),
	.c2v_87_in2 (c2v_out2[87]),
	.ch_msg_88 (ch_msg_88[DATAPATH_WIDTH-1:0]),
	.c2v_88_in0 (c2v_out0[88]),
	.c2v_88_in1 (c2v_out1[88]),
	.c2v_88_in2 (c2v_out2[88]),
	.ch_msg_89 (ch_msg_89[DATAPATH_WIDTH-1:0]),
	.c2v_89_in0 (c2v_out0[89]),
	.c2v_89_in1 (c2v_out1[89]),
	.c2v_89_in2 (c2v_out2[89]),
	.ch_msg_90 (ch_msg_90[DATAPATH_WIDTH-1:0]),
	.c2v_90_in0 (c2v_out0[90]),
	.c2v_90_in1 (c2v_out1[90]),
	.c2v_90_in2 (c2v_out2[90]),
	.ch_msg_91 (ch_msg_91[DATAPATH_WIDTH-1:0]),
	.c2v_91_in0 (c2v_out0[91]),
	.c2v_91_in1 (c2v_out1[91]),
	.c2v_91_in2 (c2v_out2[91]),
	.ch_msg_92 (ch_msg_92[DATAPATH_WIDTH-1:0]),
	.c2v_92_in0 (c2v_out0[92]),
	.c2v_92_in1 (c2v_out1[92]),
	.c2v_92_in2 (c2v_out2[92]),
	.ch_msg_93 (ch_msg_93[DATAPATH_WIDTH-1:0]),
	.c2v_93_in0 (c2v_out0[93]),
	.c2v_93_in1 (c2v_out1[93]),
	.c2v_93_in2 (c2v_out2[93]),
	.ch_msg_94 (ch_msg_94[DATAPATH_WIDTH-1:0]),
	.c2v_94_in0 (c2v_out0[94]),
	.c2v_94_in1 (c2v_out1[94]),
	.c2v_94_in2 (c2v_out2[94]),
	.ch_msg_95 (ch_msg_95[DATAPATH_WIDTH-1:0]),
	.c2v_95_in0 (c2v_out0[95]),
	.c2v_95_in1 (c2v_out1[95]),
	.c2v_95_in2 (c2v_out2[95]),
	.ch_msg_96 (ch_msg_96[DATAPATH_WIDTH-1:0]),
	.c2v_96_in0 (c2v_out0[96]),
	.c2v_96_in1 (c2v_out1[96]),
	.c2v_96_in2 (c2v_out2[96]),
	.ch_msg_97 (ch_msg_97[DATAPATH_WIDTH-1:0]),
	.c2v_97_in0 (c2v_out0[97]),
	.c2v_97_in1 (c2v_out1[97]),
	.c2v_97_in2 (c2v_out2[97]),
	.ch_msg_98 (ch_msg_98[DATAPATH_WIDTH-1:0]),
	.c2v_98_in0 (c2v_out0[98]),
	.c2v_98_in1 (c2v_out1[98]),
	.c2v_98_in2 (c2v_out2[98]),
	.ch_msg_99 (ch_msg_99[DATAPATH_WIDTH-1:0]),
	.c2v_99_in0 (c2v_out0[99]),
	.c2v_99_in1 (c2v_out1[99]),
	.c2v_99_in2 (c2v_out2[99]),
	.ch_msg_100 (ch_msg_100[DATAPATH_WIDTH-1:0]),
	.c2v_100_in0 (c2v_out0[100]),
	.c2v_100_in1 (c2v_out1[100]),
	.c2v_100_in2 (c2v_out2[100]),
	.ch_msg_101 (ch_msg_101[DATAPATH_WIDTH-1:0]),
	.c2v_101_in0 (c2v_out0[101]),
	.c2v_101_in1 (c2v_out1[101]),
	.c2v_101_in2 (c2v_out2[101]),
	.ch_msg_102 (ch_msg_102[DATAPATH_WIDTH-1:0]),
	.c2v_102_in0 (c2v_out0[102]),
	.c2v_102_in1 (c2v_out1[102]),
	.c2v_102_in2 (c2v_out2[102]),
	.ch_msg_103 (ch_msg_103[DATAPATH_WIDTH-1:0]),
	.c2v_103_in0 (c2v_out0[103]),
	.c2v_103_in1 (c2v_out1[103]),
	.c2v_103_in2 (c2v_out2[103]),
	.ch_msg_104 (ch_msg_104[DATAPATH_WIDTH-1:0]),
	.c2v_104_in0 (c2v_out0[104]),
	.c2v_104_in1 (c2v_out1[104]),
	.c2v_104_in2 (c2v_out2[104]),
	.ch_msg_105 (ch_msg_105[DATAPATH_WIDTH-1:0]),
	.c2v_105_in0 (c2v_out0[105]),
	.c2v_105_in1 (c2v_out1[105]),
	.c2v_105_in2 (c2v_out2[105]),
	.ch_msg_106 (ch_msg_106[DATAPATH_WIDTH-1:0]),
	.c2v_106_in0 (c2v_out0[106]),
	.c2v_106_in1 (c2v_out1[106]),
	.c2v_106_in2 (c2v_out2[106]),
	.ch_msg_107 (ch_msg_107[DATAPATH_WIDTH-1:0]),
	.c2v_107_in0 (c2v_out0[107]),
	.c2v_107_in1 (c2v_out1[107]),
	.c2v_107_in2 (c2v_out2[107]),
	.ch_msg_108 (ch_msg_108[DATAPATH_WIDTH-1:0]),
	.c2v_108_in0 (c2v_out0[108]),
	.c2v_108_in1 (c2v_out1[108]),
	.c2v_108_in2 (c2v_out2[108]),
	.ch_msg_109 (ch_msg_109[DATAPATH_WIDTH-1:0]),
	.c2v_109_in0 (c2v_out0[109]),
	.c2v_109_in1 (c2v_out1[109]),
	.c2v_109_in2 (c2v_out2[109]),
	.ch_msg_110 (ch_msg_110[DATAPATH_WIDTH-1:0]),
	.c2v_110_in0 (c2v_out0[110]),
	.c2v_110_in1 (c2v_out1[110]),
	.c2v_110_in2 (c2v_out2[110]),
	.ch_msg_111 (ch_msg_111[DATAPATH_WIDTH-1:0]),
	.c2v_111_in0 (c2v_out0[111]),
	.c2v_111_in1 (c2v_out1[111]),
	.c2v_111_in2 (c2v_out2[111]),
	.ch_msg_112 (ch_msg_112[DATAPATH_WIDTH-1:0]),
	.c2v_112_in0 (c2v_out0[112]),
	.c2v_112_in1 (c2v_out1[112]),
	.c2v_112_in2 (c2v_out2[112]),
	.ch_msg_113 (ch_msg_113[DATAPATH_WIDTH-1:0]),
	.c2v_113_in0 (c2v_out0[113]),
	.c2v_113_in1 (c2v_out1[113]),
	.c2v_113_in2 (c2v_out2[113]),
	.ch_msg_114 (ch_msg_114[DATAPATH_WIDTH-1:0]),
	.c2v_114_in0 (c2v_out0[114]),
	.c2v_114_in1 (c2v_out1[114]),
	.c2v_114_in2 (c2v_out2[114]),
	.ch_msg_115 (ch_msg_115[DATAPATH_WIDTH-1:0]),
	.c2v_115_in0 (c2v_out0[115]),
	.c2v_115_in1 (c2v_out1[115]),
	.c2v_115_in2 (c2v_out2[115]),
	.ch_msg_116 (ch_msg_116[DATAPATH_WIDTH-1:0]),
	.c2v_116_in0 (c2v_out0[116]),
	.c2v_116_in1 (c2v_out1[116]),
	.c2v_116_in2 (c2v_out2[116]),
	.ch_msg_117 (ch_msg_117[DATAPATH_WIDTH-1:0]),
	.c2v_117_in0 (c2v_out0[117]),
	.c2v_117_in1 (c2v_out1[117]),
	.c2v_117_in2 (c2v_out2[117]),
	.ch_msg_118 (ch_msg_118[DATAPATH_WIDTH-1:0]),
	.c2v_118_in0 (c2v_out0[118]),
	.c2v_118_in1 (c2v_out1[118]),
	.c2v_118_in2 (c2v_out2[118]),
	.ch_msg_119 (ch_msg_119[DATAPATH_WIDTH-1:0]),
	.c2v_119_in0 (c2v_out0[119]),
	.c2v_119_in1 (c2v_out1[119]),
	.c2v_119_in2 (c2v_out2[119]),
	.ch_msg_120 (ch_msg_120[DATAPATH_WIDTH-1:0]),
	.c2v_120_in0 (c2v_out0[120]),
	.c2v_120_in1 (c2v_out1[120]),
	.c2v_120_in2 (c2v_out2[120]),
	.ch_msg_121 (ch_msg_121[DATAPATH_WIDTH-1:0]),
	.c2v_121_in0 (c2v_out0[121]),
	.c2v_121_in1 (c2v_out1[121]),
	.c2v_121_in2 (c2v_out2[121]),
	.ch_msg_122 (ch_msg_122[DATAPATH_WIDTH-1:0]),
	.c2v_122_in0 (c2v_out0[122]),
	.c2v_122_in1 (c2v_out1[122]),
	.c2v_122_in2 (c2v_out2[122]),
	.ch_msg_123 (ch_msg_123[DATAPATH_WIDTH-1:0]),
	.c2v_123_in0 (c2v_out0[123]),
	.c2v_123_in1 (c2v_out1[123]),
	.c2v_123_in2 (c2v_out2[123]),
	.ch_msg_124 (ch_msg_124[DATAPATH_WIDTH-1:0]),
	.c2v_124_in0 (c2v_out0[124]),
	.c2v_124_in1 (c2v_out1[124]),
	.c2v_124_in2 (c2v_out2[124]),
	.ch_msg_125 (ch_msg_125[DATAPATH_WIDTH-1:0]),
	.c2v_125_in0 (c2v_out0[125]),
	.c2v_125_in1 (c2v_out1[125]),
	.c2v_125_in2 (c2v_out2[125]),
	.ch_msg_126 (ch_msg_126[DATAPATH_WIDTH-1:0]),
	.c2v_126_in0 (c2v_out0[126]),
	.c2v_126_in1 (c2v_out1[126]),
	.c2v_126_in2 (c2v_out2[126]),
	.ch_msg_127 (ch_msg_127[DATAPATH_WIDTH-1:0]),
	.c2v_127_in0 (c2v_out0[127]),
	.c2v_127_in1 (c2v_out1[127]),
	.c2v_127_in2 (c2v_out2[127]),
	.ch_msg_128 (ch_msg_128[DATAPATH_WIDTH-1:0]),
	.c2v_128_in0 (c2v_out0[128]),
	.c2v_128_in1 (c2v_out1[128]),
	.c2v_128_in2 (c2v_out2[128]),
	.ch_msg_129 (ch_msg_129[DATAPATH_WIDTH-1:0]),
	.c2v_129_in0 (c2v_out0[129]),
	.c2v_129_in1 (c2v_out1[129]),
	.c2v_129_in2 (c2v_out2[129]),
	.ch_msg_130 (ch_msg_130[DATAPATH_WIDTH-1:0]),
	.c2v_130_in0 (c2v_out0[130]),
	.c2v_130_in1 (c2v_out1[130]),
	.c2v_130_in2 (c2v_out2[130]),
	.ch_msg_131 (ch_msg_131[DATAPATH_WIDTH-1:0]),
	.c2v_131_in0 (c2v_out0[131]),
	.c2v_131_in1 (c2v_out1[131]),
	.c2v_131_in2 (c2v_out2[131]),
	.ch_msg_132 (ch_msg_132[DATAPATH_WIDTH-1:0]),
	.c2v_132_in0 (c2v_out0[132]),
	.c2v_132_in1 (c2v_out1[132]),
	.c2v_132_in2 (c2v_out2[132]),
	.ch_msg_133 (ch_msg_133[DATAPATH_WIDTH-1:0]),
	.c2v_133_in0 (c2v_out0[133]),
	.c2v_133_in1 (c2v_out1[133]),
	.c2v_133_in2 (c2v_out2[133]),
	.ch_msg_134 (ch_msg_134[DATAPATH_WIDTH-1:0]),
	.c2v_134_in0 (c2v_out0[134]),
	.c2v_134_in1 (c2v_out1[134]),
	.c2v_134_in2 (c2v_out2[134]),
	.ch_msg_135 (ch_msg_135[DATAPATH_WIDTH-1:0]),
	.c2v_135_in0 (c2v_out0[135]),
	.c2v_135_in1 (c2v_out1[135]),
	.c2v_135_in2 (c2v_out2[135]),
	.ch_msg_136 (ch_msg_136[DATAPATH_WIDTH-1:0]),
	.c2v_136_in0 (c2v_out0[136]),
	.c2v_136_in1 (c2v_out1[136]),
	.c2v_136_in2 (c2v_out2[136]),
	.ch_msg_137 (ch_msg_137[DATAPATH_WIDTH-1:0]),
	.c2v_137_in0 (c2v_out0[137]),
	.c2v_137_in1 (c2v_out1[137]),
	.c2v_137_in2 (c2v_out2[137]),
	.ch_msg_138 (ch_msg_138[DATAPATH_WIDTH-1:0]),
	.c2v_138_in0 (c2v_out0[138]),
	.c2v_138_in1 (c2v_out1[138]),
	.c2v_138_in2 (c2v_out2[138]),
	.ch_msg_139 (ch_msg_139[DATAPATH_WIDTH-1:0]),
	.c2v_139_in0 (c2v_out0[139]),
	.c2v_139_in1 (c2v_out1[139]),
	.c2v_139_in2 (c2v_out2[139]),
	.ch_msg_140 (ch_msg_140[DATAPATH_WIDTH-1:0]),
	.c2v_140_in0 (c2v_out0[140]),
	.c2v_140_in1 (c2v_out1[140]),
	.c2v_140_in2 (c2v_out2[140]),
	.ch_msg_141 (ch_msg_141[DATAPATH_WIDTH-1:0]),
	.c2v_141_in0 (c2v_out0[141]),
	.c2v_141_in1 (c2v_out1[141]),
	.c2v_141_in2 (c2v_out2[141]),
	.ch_msg_142 (ch_msg_142[DATAPATH_WIDTH-1:0]),
	.c2v_142_in0 (c2v_out0[142]),
	.c2v_142_in1 (c2v_out1[142]),
	.c2v_142_in2 (c2v_out2[142]),
	.ch_msg_143 (ch_msg_143[DATAPATH_WIDTH-1:0]),
	.c2v_143_in0 (c2v_out0[143]),
	.c2v_143_in1 (c2v_out1[143]),
	.c2v_143_in2 (c2v_out2[143]),
	.ch_msg_144 (ch_msg_144[DATAPATH_WIDTH-1:0]),
	.c2v_144_in0 (c2v_out0[144]),
	.c2v_144_in1 (c2v_out1[144]),
	.c2v_144_in2 (c2v_out2[144]),
	.ch_msg_145 (ch_msg_145[DATAPATH_WIDTH-1:0]),
	.c2v_145_in0 (c2v_out0[145]),
	.c2v_145_in1 (c2v_out1[145]),
	.c2v_145_in2 (c2v_out2[145]),
	.ch_msg_146 (ch_msg_146[DATAPATH_WIDTH-1:0]),
	.c2v_146_in0 (c2v_out0[146]),
	.c2v_146_in1 (c2v_out1[146]),
	.c2v_146_in2 (c2v_out2[146]),
	.ch_msg_147 (ch_msg_147[DATAPATH_WIDTH-1:0]),
	.c2v_147_in0 (c2v_out0[147]),
	.c2v_147_in1 (c2v_out1[147]),
	.c2v_147_in2 (c2v_out2[147]),
	.ch_msg_148 (ch_msg_148[DATAPATH_WIDTH-1:0]),
	.c2v_148_in0 (c2v_out0[148]),
	.c2v_148_in1 (c2v_out1[148]),
	.c2v_148_in2 (c2v_out2[148]),
	.ch_msg_149 (ch_msg_149[DATAPATH_WIDTH-1:0]),
	.c2v_149_in0 (c2v_out0[149]),
	.c2v_149_in1 (c2v_out1[149]),
	.c2v_149_in2 (c2v_out2[149]),
	.ch_msg_150 (ch_msg_150[DATAPATH_WIDTH-1:0]),
	.c2v_150_in0 (c2v_out0[150]),
	.c2v_150_in1 (c2v_out1[150]),
	.c2v_150_in2 (c2v_out2[150]),
	.ch_msg_151 (ch_msg_151[DATAPATH_WIDTH-1:0]),
	.c2v_151_in0 (c2v_out0[151]),
	.c2v_151_in1 (c2v_out1[151]),
	.c2v_151_in2 (c2v_out2[151]),
	.ch_msg_152 (ch_msg_152[DATAPATH_WIDTH-1:0]),
	.c2v_152_in0 (c2v_out0[152]),
	.c2v_152_in1 (c2v_out1[152]),
	.c2v_152_in2 (c2v_out2[152]),
	.ch_msg_153 (ch_msg_153[DATAPATH_WIDTH-1:0]),
	.c2v_153_in0 (c2v_out0[153]),
	.c2v_153_in1 (c2v_out1[153]),
	.c2v_153_in2 (c2v_out2[153]),
	.ch_msg_154 (ch_msg_154[DATAPATH_WIDTH-1:0]),
	.c2v_154_in0 (c2v_out0[154]),
	.c2v_154_in1 (c2v_out1[154]),
	.c2v_154_in2 (c2v_out2[154]),
	.ch_msg_155 (ch_msg_155[DATAPATH_WIDTH-1:0]),
	.c2v_155_in0 (c2v_out0[155]),
	.c2v_155_in1 (c2v_out1[155]),
	.c2v_155_in2 (c2v_out2[155]),
	.ch_msg_156 (ch_msg_156[DATAPATH_WIDTH-1:0]),
	.c2v_156_in0 (c2v_out0[156]),
	.c2v_156_in1 (c2v_out1[156]),
	.c2v_156_in2 (c2v_out2[156]),
	.ch_msg_157 (ch_msg_157[DATAPATH_WIDTH-1:0]),
	.c2v_157_in0 (c2v_out0[157]),
	.c2v_157_in1 (c2v_out1[157]),
	.c2v_157_in2 (c2v_out2[157]),
	.ch_msg_158 (ch_msg_158[DATAPATH_WIDTH-1:0]),
	.c2v_158_in0 (c2v_out0[158]),
	.c2v_158_in1 (c2v_out1[158]),
	.c2v_158_in2 (c2v_out2[158]),
	.ch_msg_159 (ch_msg_159[DATAPATH_WIDTH-1:0]),
	.c2v_159_in0 (c2v_out0[159]),
	.c2v_159_in1 (c2v_out1[159]),
	.c2v_159_in2 (c2v_out2[159]),
	.ch_msg_160 (ch_msg_160[DATAPATH_WIDTH-1:0]),
	.c2v_160_in0 (c2v_out0[160]),
	.c2v_160_in1 (c2v_out1[160]),
	.c2v_160_in2 (c2v_out2[160]),
	.ch_msg_161 (ch_msg_161[DATAPATH_WIDTH-1:0]),
	.c2v_161_in0 (c2v_out0[161]),
	.c2v_161_in1 (c2v_out1[161]),
	.c2v_161_in2 (c2v_out2[161]),
	.ch_msg_162 (ch_msg_162[DATAPATH_WIDTH-1:0]),
	.c2v_162_in0 (c2v_out0[162]),
	.c2v_162_in1 (c2v_out1[162]),
	.c2v_162_in2 (c2v_out2[162]),
	.ch_msg_163 (ch_msg_163[DATAPATH_WIDTH-1:0]),
	.c2v_163_in0 (c2v_out0[163]),
	.c2v_163_in1 (c2v_out1[163]),
	.c2v_163_in2 (c2v_out2[163]),
	.ch_msg_164 (ch_msg_164[DATAPATH_WIDTH-1:0]),
	.c2v_164_in0 (c2v_out0[164]),
	.c2v_164_in1 (c2v_out1[164]),
	.c2v_164_in2 (c2v_out2[164]),
	.ch_msg_165 (ch_msg_165[DATAPATH_WIDTH-1:0]),
	.c2v_165_in0 (c2v_out0[165]),
	.c2v_165_in1 (c2v_out1[165]),
	.c2v_165_in2 (c2v_out2[165]),
	.ch_msg_166 (ch_msg_166[DATAPATH_WIDTH-1:0]),
	.c2v_166_in0 (c2v_out0[166]),
	.c2v_166_in1 (c2v_out1[166]),
	.c2v_166_in2 (c2v_out2[166]),
	.ch_msg_167 (ch_msg_167[DATAPATH_WIDTH-1:0]),
	.c2v_167_in0 (c2v_out0[167]),
	.c2v_167_in1 (c2v_out1[167]),
	.c2v_167_in2 (c2v_out2[167]),
	.ch_msg_168 (ch_msg_168[DATAPATH_WIDTH-1:0]),
	.c2v_168_in0 (c2v_out0[168]),
	.c2v_168_in1 (c2v_out1[168]),
	.c2v_168_in2 (c2v_out2[168]),
	.ch_msg_169 (ch_msg_169[DATAPATH_WIDTH-1:0]),
	.c2v_169_in0 (c2v_out0[169]),
	.c2v_169_in1 (c2v_out1[169]),
	.c2v_169_in2 (c2v_out2[169]),
	.ch_msg_170 (ch_msg_170[DATAPATH_WIDTH-1:0]),
	.c2v_170_in0 (c2v_out0[170]),
	.c2v_170_in1 (c2v_out1[170]),
	.c2v_170_in2 (c2v_out2[170]),
	.ch_msg_171 (ch_msg_171[DATAPATH_WIDTH-1:0]),
	.c2v_171_in0 (c2v_out0[171]),
	.c2v_171_in1 (c2v_out1[171]),
	.c2v_171_in2 (c2v_out2[171]),
	.ch_msg_172 (ch_msg_172[DATAPATH_WIDTH-1:0]),
	.c2v_172_in0 (c2v_out0[172]),
	.c2v_172_in1 (c2v_out1[172]),
	.c2v_172_in2 (c2v_out2[172]),
	.ch_msg_173 (ch_msg_173[DATAPATH_WIDTH-1:0]),
	.c2v_173_in0 (c2v_out0[173]),
	.c2v_173_in1 (c2v_out1[173]),
	.c2v_173_in2 (c2v_out2[173]),
	.ch_msg_174 (ch_msg_174[DATAPATH_WIDTH-1:0]),
	.c2v_174_in0 (c2v_out0[174]),
	.c2v_174_in1 (c2v_out1[174]),
	.c2v_174_in2 (c2v_out2[174]),
	.ch_msg_175 (ch_msg_175[DATAPATH_WIDTH-1:0]),
	.c2v_175_in0 (c2v_out0[175]),
	.c2v_175_in1 (c2v_out1[175]),
	.c2v_175_in2 (c2v_out2[175]),
	.ch_msg_176 (ch_msg_176[DATAPATH_WIDTH-1:0]),
	.c2v_176_in0 (c2v_out0[176]),
	.c2v_176_in1 (c2v_out1[176]),
	.c2v_176_in2 (c2v_out2[176]),
	.ch_msg_177 (ch_msg_177[DATAPATH_WIDTH-1:0]),
	.c2v_177_in0 (c2v_out0[177]),
	.c2v_177_in1 (c2v_out1[177]),
	.c2v_177_in2 (c2v_out2[177]),
	.ch_msg_178 (ch_msg_178[DATAPATH_WIDTH-1:0]),
	.c2v_178_in0 (c2v_out0[178]),
	.c2v_178_in1 (c2v_out1[178]),
	.c2v_178_in2 (c2v_out2[178]),
	.ch_msg_179 (ch_msg_179[DATAPATH_WIDTH-1:0]),
	.c2v_179_in0 (c2v_out0[179]),
	.c2v_179_in1 (c2v_out1[179]),
	.c2v_179_in2 (c2v_out2[179]),
	.ch_msg_180 (ch_msg_180[DATAPATH_WIDTH-1:0]),
	.c2v_180_in0 (c2v_out0[180]),
	.c2v_180_in1 (c2v_out1[180]),
	.c2v_180_in2 (c2v_out2[180]),
	.ch_msg_181 (ch_msg_181[DATAPATH_WIDTH-1:0]),
	.c2v_181_in0 (c2v_out0[181]),
	.c2v_181_in1 (c2v_out1[181]),
	.c2v_181_in2 (c2v_out2[181]),
	.ch_msg_182 (ch_msg_182[DATAPATH_WIDTH-1:0]),
	.c2v_182_in0 (c2v_out0[182]),
	.c2v_182_in1 (c2v_out1[182]),
	.c2v_182_in2 (c2v_out2[182]),
	.ch_msg_183 (ch_msg_183[DATAPATH_WIDTH-1:0]),
	.c2v_183_in0 (c2v_out0[183]),
	.c2v_183_in1 (c2v_out1[183]),
	.c2v_183_in2 (c2v_out2[183]),
	.ch_msg_184 (ch_msg_184[DATAPATH_WIDTH-1:0]),
	.c2v_184_in0 (c2v_out0[184]),
	.c2v_184_in1 (c2v_out1[184]),
	.c2v_184_in2 (c2v_out2[184]),
	.ch_msg_185 (ch_msg_185[DATAPATH_WIDTH-1:0]),
	.c2v_185_in0 (c2v_out0[185]),
	.c2v_185_in1 (c2v_out1[185]),
	.c2v_185_in2 (c2v_out2[185]),
	.ch_msg_186 (ch_msg_186[DATAPATH_WIDTH-1:0]),
	.c2v_186_in0 (c2v_out0[186]),
	.c2v_186_in1 (c2v_out1[186]),
	.c2v_186_in2 (c2v_out2[186]),
	.ch_msg_187 (ch_msg_187[DATAPATH_WIDTH-1:0]),
	.c2v_187_in0 (c2v_out0[187]),
	.c2v_187_in1 (c2v_out1[187]),
	.c2v_187_in2 (c2v_out2[187]),
	.ch_msg_188 (ch_msg_188[DATAPATH_WIDTH-1:0]),
	.c2v_188_in0 (c2v_out0[188]),
	.c2v_188_in1 (c2v_out1[188]),
	.c2v_188_in2 (c2v_out2[188]),
	.ch_msg_189 (ch_msg_189[DATAPATH_WIDTH-1:0]),
	.c2v_189_in0 (c2v_out0[189]),
	.c2v_189_in1 (c2v_out1[189]),
	.c2v_189_in2 (c2v_out2[189]),
	.ch_msg_190 (ch_msg_190[DATAPATH_WIDTH-1:0]),
	.c2v_190_in0 (c2v_out0[190]),
	.c2v_190_in1 (c2v_out1[190]),
	.c2v_190_in2 (c2v_out2[190]),
	.ch_msg_191 (ch_msg_191[DATAPATH_WIDTH-1:0]),
	.c2v_191_in0 (c2v_out0[191]),
	.c2v_191_in1 (c2v_out1[191]),
	.c2v_191_in2 (c2v_out2[191]),
	.ch_msg_192 (ch_msg_192[DATAPATH_WIDTH-1:0]),
	.c2v_192_in0 (c2v_out0[192]),
	.c2v_192_in1 (c2v_out1[192]),
	.c2v_192_in2 (c2v_out2[192]),
	.ch_msg_193 (ch_msg_193[DATAPATH_WIDTH-1:0]),
	.c2v_193_in0 (c2v_out0[193]),
	.c2v_193_in1 (c2v_out1[193]),
	.c2v_193_in2 (c2v_out2[193]),
	.ch_msg_194 (ch_msg_194[DATAPATH_WIDTH-1:0]),
	.c2v_194_in0 (c2v_out0[194]),
	.c2v_194_in1 (c2v_out1[194]),
	.c2v_194_in2 (c2v_out2[194]),
	.ch_msg_195 (ch_msg_195[DATAPATH_WIDTH-1:0]),
	.c2v_195_in0 (c2v_out0[195]),
	.c2v_195_in1 (c2v_out1[195]),
	.c2v_195_in2 (c2v_out2[195]),
	.ch_msg_196 (ch_msg_196[DATAPATH_WIDTH-1:0]),
	.c2v_196_in0 (c2v_out0[196]),
	.c2v_196_in1 (c2v_out1[196]),
	.c2v_196_in2 (c2v_out2[196]),
	.ch_msg_197 (ch_msg_197[DATAPATH_WIDTH-1:0]),
	.c2v_197_in0 (c2v_out0[197]),
	.c2v_197_in1 (c2v_out1[197]),
	.c2v_197_in2 (c2v_out2[197]),
	.ch_msg_198 (ch_msg_198[DATAPATH_WIDTH-1:0]),
	.c2v_198_in0 (c2v_out0[198]),
	.c2v_198_in1 (c2v_out1[198]),
	.c2v_198_in2 (c2v_out2[198]),
	.ch_msg_199 (ch_msg_199[DATAPATH_WIDTH-1:0]),
	.c2v_199_in0 (c2v_out0[199]),
	.c2v_199_in1 (c2v_out1[199]),
	.c2v_199_in2 (c2v_out2[199]),
	.ch_msg_200 (ch_msg_200[DATAPATH_WIDTH-1:0]),
	.c2v_200_in0 (c2v_out0[200]),
	.c2v_200_in1 (c2v_out1[200]),
	.c2v_200_in2 (c2v_out2[200]),
	.ch_msg_201 (ch_msg_201[DATAPATH_WIDTH-1:0]),
	.c2v_201_in0 (c2v_out0[201]),
	.c2v_201_in1 (c2v_out1[201]),
	.c2v_201_in2 (c2v_out2[201]),
	.ch_msg_202 (ch_msg_202[DATAPATH_WIDTH-1:0]),
	.c2v_202_in0 (c2v_out0[202]),
	.c2v_202_in1 (c2v_out1[202]),
	.c2v_202_in2 (c2v_out2[202]),
	.ch_msg_203 (ch_msg_203[DATAPATH_WIDTH-1:0]),
	.c2v_203_in0 (c2v_out0[203]),
	.c2v_203_in1 (c2v_out1[203]),
	.c2v_203_in2 (c2v_out2[203]),

	.read_clk (read_clk),
	.read_addr_offset (vnu_read_addr_offset),
	.v2c_src (v2c_src),
	.c2v_latch_en (c2v_latch_en),
	.c2v_parallel_load (load[0]),

	// Iteration-Refresh Page Address
	.page_addr_ram_0 (vnu_page_addr_ram_0[VN_PAGE_ADDR_BW+1-1:0]),
	.page_addr_ram_1 (vnu_page_addr_ram_1[VN_PAGE_ADDR_BW+1-1:0]),
	.page_addr_ram_2 (vnu_page_addr_ram_2[DN_PAGE_ADDR_BW+1-1:0]), // the last one is for decision node
	//Iteration-Refresh Page Data
	.ram_write_dataA_0 (vnu_ram_write_dataA_0[VN_ROM_RD_BW-1:0]), // from portA of IB-ROM
	.ram_write_dataB_0 (vnu_ram_write_dataB_0[VN_ROM_RD_BW-1:0]), // from portB of IB-ROM
	.ram_write_dataA_1 (vnu_ram_write_dataA_1[VN_ROM_RD_BW-1:0]), // from portA of IB-ROM
	.ram_write_dataB_1 (vnu_ram_write_dataB_1[VN_ROM_RD_BW-1:0]), // from portB of IB-ROM
	.ram_write_dataA_2 (vnu_ram_write_dataA_2[DN_ROM_RD_BW-1:0]), // from portA of IB-ROM (for decision node)
	.ram_write_dataB_2 (vnu_ram_write_dataB_2[DN_ROM_RD_BW-1:0]), // from portB of IB-ROM (for decision node)
	.ib_ram_we (vnu_ib_ram_we[IB_VNU_DECOMP_funNum:0]),
	.vn_write_clk (vn_write_clk),
	.dn_write_clk (dn_write_clk)
);


 // Instatiation of Routing Network and Port Mapping
fully_parallel_route #(
	.DATAPATH_WIDTH(DATAPATH_WIDTH),
	.CN_DEGREE     (CN_DEGREE),
	.VN_DEGREE     (VN_DEGREE),
	.MSG_WIDTH     (MSG_WIDTH)
) routing_network (
// (N-K) number of check-to-Variable message buses, each of which is d_c bit width as input ports of this routing network
	.v2c_parallelOut_00(v2c_out0[0]),
	.v2c_parallelOut_01(v2c_out1[0]),
	.v2c_parallelOut_02(v2c_out2[0]),
	.v2c_parallelOut_03(v2c_out3[0]),
	.v2c_parallelOut_04(v2c_out4[0]),
	.v2c_parallelOut_05(v2c_out5[0]),
	.v2c_parallelOut_10(v2c_out0[1]),
	.v2c_parallelOut_11(v2c_out1[1]),
	.v2c_parallelOut_12(v2c_out2[1]),
	.v2c_parallelOut_13(v2c_out3[1]),
	.v2c_parallelOut_14(v2c_out4[1]),
	.v2c_parallelOut_15(v2c_out5[1]),
	.v2c_parallelOut_20(v2c_out0[2]),
	.v2c_parallelOut_21(v2c_out1[2]),
	.v2c_parallelOut_22(v2c_out2[2]),
	.v2c_parallelOut_23(v2c_out3[2]),
	.v2c_parallelOut_24(v2c_out4[2]),
	.v2c_parallelOut_25(v2c_out5[2]),
	.v2c_parallelOut_30(v2c_out0[3]),
	.v2c_parallelOut_31(v2c_out1[3]),
	.v2c_parallelOut_32(v2c_out2[3]),
	.v2c_parallelOut_33(v2c_out3[3]),
	.v2c_parallelOut_34(v2c_out4[3]),
	.v2c_parallelOut_35(v2c_out5[3]),
	.v2c_parallelOut_40(v2c_out0[4]),
	.v2c_parallelOut_41(v2c_out1[4]),
	.v2c_parallelOut_42(v2c_out2[4]),
	.v2c_parallelOut_43(v2c_out3[4]),
	.v2c_parallelOut_44(v2c_out4[4]),
	.v2c_parallelOut_45(v2c_out5[4]),
	.v2c_parallelOut_50(v2c_out0[5]),
	.v2c_parallelOut_51(v2c_out1[5]),
	.v2c_parallelOut_52(v2c_out2[5]),
	.v2c_parallelOut_53(v2c_out3[5]),
	.v2c_parallelOut_54(v2c_out4[5]),
	.v2c_parallelOut_55(v2c_out5[5]),
	.v2c_parallelOut_60(v2c_out0[6]),
	.v2c_parallelOut_61(v2c_out1[6]),
	.v2c_parallelOut_62(v2c_out2[6]),
	.v2c_parallelOut_63(v2c_out3[6]),
	.v2c_parallelOut_64(v2c_out4[6]),
	.v2c_parallelOut_65(v2c_out5[6]),
	.v2c_parallelOut_70(v2c_out0[7]),
	.v2c_parallelOut_71(v2c_out1[7]),
	.v2c_parallelOut_72(v2c_out2[7]),
	.v2c_parallelOut_73(v2c_out3[7]),
	.v2c_parallelOut_74(v2c_out4[7]),
	.v2c_parallelOut_75(v2c_out5[7]),
	.v2c_parallelOut_80(v2c_out0[8]),
	.v2c_parallelOut_81(v2c_out1[8]),
	.v2c_parallelOut_82(v2c_out2[8]),
	.v2c_parallelOut_83(v2c_out3[8]),
	.v2c_parallelOut_84(v2c_out4[8]),
	.v2c_parallelOut_85(v2c_out5[8]),
	.v2c_parallelOut_90(v2c_out0[9]),
	.v2c_parallelOut_91(v2c_out1[9]),
	.v2c_parallelOut_92(v2c_out2[9]),
	.v2c_parallelOut_93(v2c_out3[9]),
	.v2c_parallelOut_94(v2c_out4[9]),
	.v2c_parallelOut_95(v2c_out5[9]),
	.v2c_parallelOut_100(v2c_out0[10]),
	.v2c_parallelOut_101(v2c_out1[10]),
	.v2c_parallelOut_102(v2c_out2[10]),
	.v2c_parallelOut_103(v2c_out3[10]),
	.v2c_parallelOut_104(v2c_out4[10]),
	.v2c_parallelOut_105(v2c_out5[10]),
	.v2c_parallelOut_110(v2c_out0[11]),
	.v2c_parallelOut_111(v2c_out1[11]),
	.v2c_parallelOut_112(v2c_out2[11]),
	.v2c_parallelOut_113(v2c_out3[11]),
	.v2c_parallelOut_114(v2c_out4[11]),
	.v2c_parallelOut_115(v2c_out5[11]),
	.v2c_parallelOut_120(v2c_out0[12]),
	.v2c_parallelOut_121(v2c_out1[12]),
	.v2c_parallelOut_122(v2c_out2[12]),
	.v2c_parallelOut_123(v2c_out3[12]),
	.v2c_parallelOut_124(v2c_out4[12]),
	.v2c_parallelOut_125(v2c_out5[12]),
	.v2c_parallelOut_130(v2c_out0[13]),
	.v2c_parallelOut_131(v2c_out1[13]),
	.v2c_parallelOut_132(v2c_out2[13]),
	.v2c_parallelOut_133(v2c_out3[13]),
	.v2c_parallelOut_134(v2c_out4[13]),
	.v2c_parallelOut_135(v2c_out5[13]),
	.v2c_parallelOut_140(v2c_out0[14]),
	.v2c_parallelOut_141(v2c_out1[14]),
	.v2c_parallelOut_142(v2c_out2[14]),
	.v2c_parallelOut_143(v2c_out3[14]),
	.v2c_parallelOut_144(v2c_out4[14]),
	.v2c_parallelOut_145(v2c_out5[14]),
	.v2c_parallelOut_150(v2c_out0[15]),
	.v2c_parallelOut_151(v2c_out1[15]),
	.v2c_parallelOut_152(v2c_out2[15]),
	.v2c_parallelOut_153(v2c_out3[15]),
	.v2c_parallelOut_154(v2c_out4[15]),
	.v2c_parallelOut_155(v2c_out5[15]),
	.v2c_parallelOut_160(v2c_out0[16]),
	.v2c_parallelOut_161(v2c_out1[16]),
	.v2c_parallelOut_162(v2c_out2[16]),
	.v2c_parallelOut_163(v2c_out3[16]),
	.v2c_parallelOut_164(v2c_out4[16]),
	.v2c_parallelOut_165(v2c_out5[16]),
	.v2c_parallelOut_170(v2c_out0[17]),
	.v2c_parallelOut_171(v2c_out1[17]),
	.v2c_parallelOut_172(v2c_out2[17]),
	.v2c_parallelOut_173(v2c_out3[17]),
	.v2c_parallelOut_174(v2c_out4[17]),
	.v2c_parallelOut_175(v2c_out5[17]),
	.v2c_parallelOut_180(v2c_out0[18]),
	.v2c_parallelOut_181(v2c_out1[18]),
	.v2c_parallelOut_182(v2c_out2[18]),
	.v2c_parallelOut_183(v2c_out3[18]),
	.v2c_parallelOut_184(v2c_out4[18]),
	.v2c_parallelOut_185(v2c_out5[18]),
	.v2c_parallelOut_190(v2c_out0[19]),
	.v2c_parallelOut_191(v2c_out1[19]),
	.v2c_parallelOut_192(v2c_out2[19]),
	.v2c_parallelOut_193(v2c_out3[19]),
	.v2c_parallelOut_194(v2c_out4[19]),
	.v2c_parallelOut_195(v2c_out5[19]),
	.v2c_parallelOut_200(v2c_out0[20]),
	.v2c_parallelOut_201(v2c_out1[20]),
	.v2c_parallelOut_202(v2c_out2[20]),
	.v2c_parallelOut_203(v2c_out3[20]),
	.v2c_parallelOut_204(v2c_out4[20]),
	.v2c_parallelOut_205(v2c_out5[20]),
	.v2c_parallelOut_210(v2c_out0[21]),
	.v2c_parallelOut_211(v2c_out1[21]),
	.v2c_parallelOut_212(v2c_out2[21]),
	.v2c_parallelOut_213(v2c_out3[21]),
	.v2c_parallelOut_214(v2c_out4[21]),
	.v2c_parallelOut_215(v2c_out5[21]),
	.v2c_parallelOut_220(v2c_out0[22]),
	.v2c_parallelOut_221(v2c_out1[22]),
	.v2c_parallelOut_222(v2c_out2[22]),
	.v2c_parallelOut_223(v2c_out3[22]),
	.v2c_parallelOut_224(v2c_out4[22]),
	.v2c_parallelOut_225(v2c_out5[22]),
	.v2c_parallelOut_230(v2c_out0[23]),
	.v2c_parallelOut_231(v2c_out1[23]),
	.v2c_parallelOut_232(v2c_out2[23]),
	.v2c_parallelOut_233(v2c_out3[23]),
	.v2c_parallelOut_234(v2c_out4[23]),
	.v2c_parallelOut_235(v2c_out5[23]),
	.v2c_parallelOut_240(v2c_out0[24]),
	.v2c_parallelOut_241(v2c_out1[24]),
	.v2c_parallelOut_242(v2c_out2[24]),
	.v2c_parallelOut_243(v2c_out3[24]),
	.v2c_parallelOut_244(v2c_out4[24]),
	.v2c_parallelOut_245(v2c_out5[24]),
	.v2c_parallelOut_250(v2c_out0[25]),
	.v2c_parallelOut_251(v2c_out1[25]),
	.v2c_parallelOut_252(v2c_out2[25]),
	.v2c_parallelOut_253(v2c_out3[25]),
	.v2c_parallelOut_254(v2c_out4[25]),
	.v2c_parallelOut_255(v2c_out5[25]),
	.v2c_parallelOut_260(v2c_out0[26]),
	.v2c_parallelOut_261(v2c_out1[26]),
	.v2c_parallelOut_262(v2c_out2[26]),
	.v2c_parallelOut_263(v2c_out3[26]),
	.v2c_parallelOut_264(v2c_out4[26]),
	.v2c_parallelOut_265(v2c_out5[26]),
	.v2c_parallelOut_270(v2c_out0[27]),
	.v2c_parallelOut_271(v2c_out1[27]),
	.v2c_parallelOut_272(v2c_out2[27]),
	.v2c_parallelOut_273(v2c_out3[27]),
	.v2c_parallelOut_274(v2c_out4[27]),
	.v2c_parallelOut_275(v2c_out5[27]),
	.v2c_parallelOut_280(v2c_out0[28]),
	.v2c_parallelOut_281(v2c_out1[28]),
	.v2c_parallelOut_282(v2c_out2[28]),
	.v2c_parallelOut_283(v2c_out3[28]),
	.v2c_parallelOut_284(v2c_out4[28]),
	.v2c_parallelOut_285(v2c_out5[28]),
	.v2c_parallelOut_290(v2c_out0[29]),
	.v2c_parallelOut_291(v2c_out1[29]),
	.v2c_parallelOut_292(v2c_out2[29]),
	.v2c_parallelOut_293(v2c_out3[29]),
	.v2c_parallelOut_294(v2c_out4[29]),
	.v2c_parallelOut_295(v2c_out5[29]),
	.v2c_parallelOut_300(v2c_out0[30]),
	.v2c_parallelOut_301(v2c_out1[30]),
	.v2c_parallelOut_302(v2c_out2[30]),
	.v2c_parallelOut_303(v2c_out3[30]),
	.v2c_parallelOut_304(v2c_out4[30]),
	.v2c_parallelOut_305(v2c_out5[30]),
	.v2c_parallelOut_310(v2c_out0[31]),
	.v2c_parallelOut_311(v2c_out1[31]),
	.v2c_parallelOut_312(v2c_out2[31]),
	.v2c_parallelOut_313(v2c_out3[31]),
	.v2c_parallelOut_314(v2c_out4[31]),
	.v2c_parallelOut_315(v2c_out5[31]),
	.v2c_parallelOut_320(v2c_out0[32]),
	.v2c_parallelOut_321(v2c_out1[32]),
	.v2c_parallelOut_322(v2c_out2[32]),
	.v2c_parallelOut_323(v2c_out3[32]),
	.v2c_parallelOut_324(v2c_out4[32]),
	.v2c_parallelOut_325(v2c_out5[32]),
	.v2c_parallelOut_330(v2c_out0[33]),
	.v2c_parallelOut_331(v2c_out1[33]),
	.v2c_parallelOut_332(v2c_out2[33]),
	.v2c_parallelOut_333(v2c_out3[33]),
	.v2c_parallelOut_334(v2c_out4[33]),
	.v2c_parallelOut_335(v2c_out5[33]),
	.v2c_parallelOut_340(v2c_out0[34]),
	.v2c_parallelOut_341(v2c_out1[34]),
	.v2c_parallelOut_342(v2c_out2[34]),
	.v2c_parallelOut_343(v2c_out3[34]),
	.v2c_parallelOut_344(v2c_out4[34]),
	.v2c_parallelOut_345(v2c_out5[34]),
	.v2c_parallelOut_350(v2c_out0[35]),
	.v2c_parallelOut_351(v2c_out1[35]),
	.v2c_parallelOut_352(v2c_out2[35]),
	.v2c_parallelOut_353(v2c_out3[35]),
	.v2c_parallelOut_354(v2c_out4[35]),
	.v2c_parallelOut_355(v2c_out5[35]),
	.v2c_parallelOut_360(v2c_out0[36]),
	.v2c_parallelOut_361(v2c_out1[36]),
	.v2c_parallelOut_362(v2c_out2[36]),
	.v2c_parallelOut_363(v2c_out3[36]),
	.v2c_parallelOut_364(v2c_out4[36]),
	.v2c_parallelOut_365(v2c_out5[36]),
	.v2c_parallelOut_370(v2c_out0[37]),
	.v2c_parallelOut_371(v2c_out1[37]),
	.v2c_parallelOut_372(v2c_out2[37]),
	.v2c_parallelOut_373(v2c_out3[37]),
	.v2c_parallelOut_374(v2c_out4[37]),
	.v2c_parallelOut_375(v2c_out5[37]),
	.v2c_parallelOut_380(v2c_out0[38]),
	.v2c_parallelOut_381(v2c_out1[38]),
	.v2c_parallelOut_382(v2c_out2[38]),
	.v2c_parallelOut_383(v2c_out3[38]),
	.v2c_parallelOut_384(v2c_out4[38]),
	.v2c_parallelOut_385(v2c_out5[38]),
	.v2c_parallelOut_390(v2c_out0[39]),
	.v2c_parallelOut_391(v2c_out1[39]),
	.v2c_parallelOut_392(v2c_out2[39]),
	.v2c_parallelOut_393(v2c_out3[39]),
	.v2c_parallelOut_394(v2c_out4[39]),
	.v2c_parallelOut_395(v2c_out5[39]),
	.v2c_parallelOut_400(v2c_out0[40]),
	.v2c_parallelOut_401(v2c_out1[40]),
	.v2c_parallelOut_402(v2c_out2[40]),
	.v2c_parallelOut_403(v2c_out3[40]),
	.v2c_parallelOut_404(v2c_out4[40]),
	.v2c_parallelOut_405(v2c_out5[40]),
	.v2c_parallelOut_410(v2c_out0[41]),
	.v2c_parallelOut_411(v2c_out1[41]),
	.v2c_parallelOut_412(v2c_out2[41]),
	.v2c_parallelOut_413(v2c_out3[41]),
	.v2c_parallelOut_414(v2c_out4[41]),
	.v2c_parallelOut_415(v2c_out5[41]),
	.v2c_parallelOut_420(v2c_out0[42]),
	.v2c_parallelOut_421(v2c_out1[42]),
	.v2c_parallelOut_422(v2c_out2[42]),
	.v2c_parallelOut_423(v2c_out3[42]),
	.v2c_parallelOut_424(v2c_out4[42]),
	.v2c_parallelOut_425(v2c_out5[42]),
	.v2c_parallelOut_430(v2c_out0[43]),
	.v2c_parallelOut_431(v2c_out1[43]),
	.v2c_parallelOut_432(v2c_out2[43]),
	.v2c_parallelOut_433(v2c_out3[43]),
	.v2c_parallelOut_434(v2c_out4[43]),
	.v2c_parallelOut_435(v2c_out5[43]),
	.v2c_parallelOut_440(v2c_out0[44]),
	.v2c_parallelOut_441(v2c_out1[44]),
	.v2c_parallelOut_442(v2c_out2[44]),
	.v2c_parallelOut_443(v2c_out3[44]),
	.v2c_parallelOut_444(v2c_out4[44]),
	.v2c_parallelOut_445(v2c_out5[44]),
	.v2c_parallelOut_450(v2c_out0[45]),
	.v2c_parallelOut_451(v2c_out1[45]),
	.v2c_parallelOut_452(v2c_out2[45]),
	.v2c_parallelOut_453(v2c_out3[45]),
	.v2c_parallelOut_454(v2c_out4[45]),
	.v2c_parallelOut_455(v2c_out5[45]),
	.v2c_parallelOut_460(v2c_out0[46]),
	.v2c_parallelOut_461(v2c_out1[46]),
	.v2c_parallelOut_462(v2c_out2[46]),
	.v2c_parallelOut_463(v2c_out3[46]),
	.v2c_parallelOut_464(v2c_out4[46]),
	.v2c_parallelOut_465(v2c_out5[46]),
	.v2c_parallelOut_470(v2c_out0[47]),
	.v2c_parallelOut_471(v2c_out1[47]),
	.v2c_parallelOut_472(v2c_out2[47]),
	.v2c_parallelOut_473(v2c_out3[47]),
	.v2c_parallelOut_474(v2c_out4[47]),
	.v2c_parallelOut_475(v2c_out5[47]),
	.v2c_parallelOut_480(v2c_out0[48]),
	.v2c_parallelOut_481(v2c_out1[48]),
	.v2c_parallelOut_482(v2c_out2[48]),
	.v2c_parallelOut_483(v2c_out3[48]),
	.v2c_parallelOut_484(v2c_out4[48]),
	.v2c_parallelOut_485(v2c_out5[48]),
	.v2c_parallelOut_490(v2c_out0[49]),
	.v2c_parallelOut_491(v2c_out1[49]),
	.v2c_parallelOut_492(v2c_out2[49]),
	.v2c_parallelOut_493(v2c_out3[49]),
	.v2c_parallelOut_494(v2c_out4[49]),
	.v2c_parallelOut_495(v2c_out5[49]),
	.v2c_parallelOut_500(v2c_out0[50]),
	.v2c_parallelOut_501(v2c_out1[50]),
	.v2c_parallelOut_502(v2c_out2[50]),
	.v2c_parallelOut_503(v2c_out3[50]),
	.v2c_parallelOut_504(v2c_out4[50]),
	.v2c_parallelOut_505(v2c_out5[50]),
	.v2c_parallelOut_510(v2c_out0[51]),
	.v2c_parallelOut_511(v2c_out1[51]),
	.v2c_parallelOut_512(v2c_out2[51]),
	.v2c_parallelOut_513(v2c_out3[51]),
	.v2c_parallelOut_514(v2c_out4[51]),
	.v2c_parallelOut_515(v2c_out5[51]),
	.v2c_parallelOut_520(v2c_out0[52]),
	.v2c_parallelOut_521(v2c_out1[52]),
	.v2c_parallelOut_522(v2c_out2[52]),
	.v2c_parallelOut_523(v2c_out3[52]),
	.v2c_parallelOut_524(v2c_out4[52]),
	.v2c_parallelOut_525(v2c_out5[52]),
	.v2c_parallelOut_530(v2c_out0[53]),
	.v2c_parallelOut_531(v2c_out1[53]),
	.v2c_parallelOut_532(v2c_out2[53]),
	.v2c_parallelOut_533(v2c_out3[53]),
	.v2c_parallelOut_534(v2c_out4[53]),
	.v2c_parallelOut_535(v2c_out5[53]),
	.v2c_parallelOut_540(v2c_out0[54]),
	.v2c_parallelOut_541(v2c_out1[54]),
	.v2c_parallelOut_542(v2c_out2[54]),
	.v2c_parallelOut_543(v2c_out3[54]),
	.v2c_parallelOut_544(v2c_out4[54]),
	.v2c_parallelOut_545(v2c_out5[54]),
	.v2c_parallelOut_550(v2c_out0[55]),
	.v2c_parallelOut_551(v2c_out1[55]),
	.v2c_parallelOut_552(v2c_out2[55]),
	.v2c_parallelOut_553(v2c_out3[55]),
	.v2c_parallelOut_554(v2c_out4[55]),
	.v2c_parallelOut_555(v2c_out5[55]),
	.v2c_parallelOut_560(v2c_out0[56]),
	.v2c_parallelOut_561(v2c_out1[56]),
	.v2c_parallelOut_562(v2c_out2[56]),
	.v2c_parallelOut_563(v2c_out3[56]),
	.v2c_parallelOut_564(v2c_out4[56]),
	.v2c_parallelOut_565(v2c_out5[56]),
	.v2c_parallelOut_570(v2c_out0[57]),
	.v2c_parallelOut_571(v2c_out1[57]),
	.v2c_parallelOut_572(v2c_out2[57]),
	.v2c_parallelOut_573(v2c_out3[57]),
	.v2c_parallelOut_574(v2c_out4[57]),
	.v2c_parallelOut_575(v2c_out5[57]),
	.v2c_parallelOut_580(v2c_out0[58]),
	.v2c_parallelOut_581(v2c_out1[58]),
	.v2c_parallelOut_582(v2c_out2[58]),
	.v2c_parallelOut_583(v2c_out3[58]),
	.v2c_parallelOut_584(v2c_out4[58]),
	.v2c_parallelOut_585(v2c_out5[58]),
	.v2c_parallelOut_590(v2c_out0[59]),
	.v2c_parallelOut_591(v2c_out1[59]),
	.v2c_parallelOut_592(v2c_out2[59]),
	.v2c_parallelOut_593(v2c_out3[59]),
	.v2c_parallelOut_594(v2c_out4[59]),
	.v2c_parallelOut_595(v2c_out5[59]),
	.v2c_parallelOut_600(v2c_out0[60]),
	.v2c_parallelOut_601(v2c_out1[60]),
	.v2c_parallelOut_602(v2c_out2[60]),
	.v2c_parallelOut_603(v2c_out3[60]),
	.v2c_parallelOut_604(v2c_out4[60]),
	.v2c_parallelOut_605(v2c_out5[60]),
	.v2c_parallelOut_610(v2c_out0[61]),
	.v2c_parallelOut_611(v2c_out1[61]),
	.v2c_parallelOut_612(v2c_out2[61]),
	.v2c_parallelOut_613(v2c_out3[61]),
	.v2c_parallelOut_614(v2c_out4[61]),
	.v2c_parallelOut_615(v2c_out5[61]),
	.v2c_parallelOut_620(v2c_out0[62]),
	.v2c_parallelOut_621(v2c_out1[62]),
	.v2c_parallelOut_622(v2c_out2[62]),
	.v2c_parallelOut_623(v2c_out3[62]),
	.v2c_parallelOut_624(v2c_out4[62]),
	.v2c_parallelOut_625(v2c_out5[62]),
	.v2c_parallelOut_630(v2c_out0[63]),
	.v2c_parallelOut_631(v2c_out1[63]),
	.v2c_parallelOut_632(v2c_out2[63]),
	.v2c_parallelOut_633(v2c_out3[63]),
	.v2c_parallelOut_634(v2c_out4[63]),
	.v2c_parallelOut_635(v2c_out5[63]),
	.v2c_parallelOut_640(v2c_out0[64]),
	.v2c_parallelOut_641(v2c_out1[64]),
	.v2c_parallelOut_642(v2c_out2[64]),
	.v2c_parallelOut_643(v2c_out3[64]),
	.v2c_parallelOut_644(v2c_out4[64]),
	.v2c_parallelOut_645(v2c_out5[64]),
	.v2c_parallelOut_650(v2c_out0[65]),
	.v2c_parallelOut_651(v2c_out1[65]),
	.v2c_parallelOut_652(v2c_out2[65]),
	.v2c_parallelOut_653(v2c_out3[65]),
	.v2c_parallelOut_654(v2c_out4[65]),
	.v2c_parallelOut_655(v2c_out5[65]),
	.v2c_parallelOut_660(v2c_out0[66]),
	.v2c_parallelOut_661(v2c_out1[66]),
	.v2c_parallelOut_662(v2c_out2[66]),
	.v2c_parallelOut_663(v2c_out3[66]),
	.v2c_parallelOut_664(v2c_out4[66]),
	.v2c_parallelOut_665(v2c_out5[66]),
	.v2c_parallelOut_670(v2c_out0[67]),
	.v2c_parallelOut_671(v2c_out1[67]),
	.v2c_parallelOut_672(v2c_out2[67]),
	.v2c_parallelOut_673(v2c_out3[67]),
	.v2c_parallelOut_674(v2c_out4[67]),
	.v2c_parallelOut_675(v2c_out5[67]),
	.v2c_parallelOut_680(v2c_out0[68]),
	.v2c_parallelOut_681(v2c_out1[68]),
	.v2c_parallelOut_682(v2c_out2[68]),
	.v2c_parallelOut_683(v2c_out3[68]),
	.v2c_parallelOut_684(v2c_out4[68]),
	.v2c_parallelOut_685(v2c_out5[68]),
	.v2c_parallelOut_690(v2c_out0[69]),
	.v2c_parallelOut_691(v2c_out1[69]),
	.v2c_parallelOut_692(v2c_out2[69]),
	.v2c_parallelOut_693(v2c_out3[69]),
	.v2c_parallelOut_694(v2c_out4[69]),
	.v2c_parallelOut_695(v2c_out5[69]),
	.v2c_parallelOut_700(v2c_out0[70]),
	.v2c_parallelOut_701(v2c_out1[70]),
	.v2c_parallelOut_702(v2c_out2[70]),
	.v2c_parallelOut_703(v2c_out3[70]),
	.v2c_parallelOut_704(v2c_out4[70]),
	.v2c_parallelOut_705(v2c_out5[70]),
	.v2c_parallelOut_710(v2c_out0[71]),
	.v2c_parallelOut_711(v2c_out1[71]),
	.v2c_parallelOut_712(v2c_out2[71]),
	.v2c_parallelOut_713(v2c_out3[71]),
	.v2c_parallelOut_714(v2c_out4[71]),
	.v2c_parallelOut_715(v2c_out5[71]),
	.v2c_parallelOut_720(v2c_out0[72]),
	.v2c_parallelOut_721(v2c_out1[72]),
	.v2c_parallelOut_722(v2c_out2[72]),
	.v2c_parallelOut_723(v2c_out3[72]),
	.v2c_parallelOut_724(v2c_out4[72]),
	.v2c_parallelOut_725(v2c_out5[72]),
	.v2c_parallelOut_730(v2c_out0[73]),
	.v2c_parallelOut_731(v2c_out1[73]),
	.v2c_parallelOut_732(v2c_out2[73]),
	.v2c_parallelOut_733(v2c_out3[73]),
	.v2c_parallelOut_734(v2c_out4[73]),
	.v2c_parallelOut_735(v2c_out5[73]),
	.v2c_parallelOut_740(v2c_out0[74]),
	.v2c_parallelOut_741(v2c_out1[74]),
	.v2c_parallelOut_742(v2c_out2[74]),
	.v2c_parallelOut_743(v2c_out3[74]),
	.v2c_parallelOut_744(v2c_out4[74]),
	.v2c_parallelOut_745(v2c_out5[74]),
	.v2c_parallelOut_750(v2c_out0[75]),
	.v2c_parallelOut_751(v2c_out1[75]),
	.v2c_parallelOut_752(v2c_out2[75]),
	.v2c_parallelOut_753(v2c_out3[75]),
	.v2c_parallelOut_754(v2c_out4[75]),
	.v2c_parallelOut_755(v2c_out5[75]),
	.v2c_parallelOut_760(v2c_out0[76]),
	.v2c_parallelOut_761(v2c_out1[76]),
	.v2c_parallelOut_762(v2c_out2[76]),
	.v2c_parallelOut_763(v2c_out3[76]),
	.v2c_parallelOut_764(v2c_out4[76]),
	.v2c_parallelOut_765(v2c_out5[76]),
	.v2c_parallelOut_770(v2c_out0[77]),
	.v2c_parallelOut_771(v2c_out1[77]),
	.v2c_parallelOut_772(v2c_out2[77]),
	.v2c_parallelOut_773(v2c_out3[77]),
	.v2c_parallelOut_774(v2c_out4[77]),
	.v2c_parallelOut_775(v2c_out5[77]),
	.v2c_parallelOut_780(v2c_out0[78]),
	.v2c_parallelOut_781(v2c_out1[78]),
	.v2c_parallelOut_782(v2c_out2[78]),
	.v2c_parallelOut_783(v2c_out3[78]),
	.v2c_parallelOut_784(v2c_out4[78]),
	.v2c_parallelOut_785(v2c_out5[78]),
	.v2c_parallelOut_790(v2c_out0[79]),
	.v2c_parallelOut_791(v2c_out1[79]),
	.v2c_parallelOut_792(v2c_out2[79]),
	.v2c_parallelOut_793(v2c_out3[79]),
	.v2c_parallelOut_794(v2c_out4[79]),
	.v2c_parallelOut_795(v2c_out5[79]),
	.v2c_parallelOut_800(v2c_out0[80]),
	.v2c_parallelOut_801(v2c_out1[80]),
	.v2c_parallelOut_802(v2c_out2[80]),
	.v2c_parallelOut_803(v2c_out3[80]),
	.v2c_parallelOut_804(v2c_out4[80]),
	.v2c_parallelOut_805(v2c_out5[80]),
	.v2c_parallelOut_810(v2c_out0[81]),
	.v2c_parallelOut_811(v2c_out1[81]),
	.v2c_parallelOut_812(v2c_out2[81]),
	.v2c_parallelOut_813(v2c_out3[81]),
	.v2c_parallelOut_814(v2c_out4[81]),
	.v2c_parallelOut_815(v2c_out5[81]),
	.v2c_parallelOut_820(v2c_out0[82]),
	.v2c_parallelOut_821(v2c_out1[82]),
	.v2c_parallelOut_822(v2c_out2[82]),
	.v2c_parallelOut_823(v2c_out3[82]),
	.v2c_parallelOut_824(v2c_out4[82]),
	.v2c_parallelOut_825(v2c_out5[82]),
	.v2c_parallelOut_830(v2c_out0[83]),
	.v2c_parallelOut_831(v2c_out1[83]),
	.v2c_parallelOut_832(v2c_out2[83]),
	.v2c_parallelOut_833(v2c_out3[83]),
	.v2c_parallelOut_834(v2c_out4[83]),
	.v2c_parallelOut_835(v2c_out5[83]),
	.v2c_parallelOut_840(v2c_out0[84]),
	.v2c_parallelOut_841(v2c_out1[84]),
	.v2c_parallelOut_842(v2c_out2[84]),
	.v2c_parallelOut_843(v2c_out3[84]),
	.v2c_parallelOut_844(v2c_out4[84]),
	.v2c_parallelOut_845(v2c_out5[84]),
	.v2c_parallelOut_850(v2c_out0[85]),
	.v2c_parallelOut_851(v2c_out1[85]),
	.v2c_parallelOut_852(v2c_out2[85]),
	.v2c_parallelOut_853(v2c_out3[85]),
	.v2c_parallelOut_854(v2c_out4[85]),
	.v2c_parallelOut_855(v2c_out5[85]),
	.v2c_parallelOut_860(v2c_out0[86]),
	.v2c_parallelOut_861(v2c_out1[86]),
	.v2c_parallelOut_862(v2c_out2[86]),
	.v2c_parallelOut_863(v2c_out3[86]),
	.v2c_parallelOut_864(v2c_out4[86]),
	.v2c_parallelOut_865(v2c_out5[86]),
	.v2c_parallelOut_870(v2c_out0[87]),
	.v2c_parallelOut_871(v2c_out1[87]),
	.v2c_parallelOut_872(v2c_out2[87]),
	.v2c_parallelOut_873(v2c_out3[87]),
	.v2c_parallelOut_874(v2c_out4[87]),
	.v2c_parallelOut_875(v2c_out5[87]),
	.v2c_parallelOut_880(v2c_out0[88]),
	.v2c_parallelOut_881(v2c_out1[88]),
	.v2c_parallelOut_882(v2c_out2[88]),
	.v2c_parallelOut_883(v2c_out3[88]),
	.v2c_parallelOut_884(v2c_out4[88]),
	.v2c_parallelOut_885(v2c_out5[88]),
	.v2c_parallelOut_890(v2c_out0[89]),
	.v2c_parallelOut_891(v2c_out1[89]),
	.v2c_parallelOut_892(v2c_out2[89]),
	.v2c_parallelOut_893(v2c_out3[89]),
	.v2c_parallelOut_894(v2c_out4[89]),
	.v2c_parallelOut_895(v2c_out5[89]),
	.v2c_parallelOut_900(v2c_out0[90]),
	.v2c_parallelOut_901(v2c_out1[90]),
	.v2c_parallelOut_902(v2c_out2[90]),
	.v2c_parallelOut_903(v2c_out3[90]),
	.v2c_parallelOut_904(v2c_out4[90]),
	.v2c_parallelOut_905(v2c_out5[90]),
	.v2c_parallelOut_910(v2c_out0[91]),
	.v2c_parallelOut_911(v2c_out1[91]),
	.v2c_parallelOut_912(v2c_out2[91]),
	.v2c_parallelOut_913(v2c_out3[91]),
	.v2c_parallelOut_914(v2c_out4[91]),
	.v2c_parallelOut_915(v2c_out5[91]),
	.v2c_parallelOut_920(v2c_out0[92]),
	.v2c_parallelOut_921(v2c_out1[92]),
	.v2c_parallelOut_922(v2c_out2[92]),
	.v2c_parallelOut_923(v2c_out3[92]),
	.v2c_parallelOut_924(v2c_out4[92]),
	.v2c_parallelOut_925(v2c_out5[92]),
	.v2c_parallelOut_930(v2c_out0[93]),
	.v2c_parallelOut_931(v2c_out1[93]),
	.v2c_parallelOut_932(v2c_out2[93]),
	.v2c_parallelOut_933(v2c_out3[93]),
	.v2c_parallelOut_934(v2c_out4[93]),
	.v2c_parallelOut_935(v2c_out5[93]),
	.v2c_parallelOut_940(v2c_out0[94]),
	.v2c_parallelOut_941(v2c_out1[94]),
	.v2c_parallelOut_942(v2c_out2[94]),
	.v2c_parallelOut_943(v2c_out3[94]),
	.v2c_parallelOut_944(v2c_out4[94]),
	.v2c_parallelOut_945(v2c_out5[94]),
	.v2c_parallelOut_950(v2c_out0[95]),
	.v2c_parallelOut_951(v2c_out1[95]),
	.v2c_parallelOut_952(v2c_out2[95]),
	.v2c_parallelOut_953(v2c_out3[95]),
	.v2c_parallelOut_954(v2c_out4[95]),
	.v2c_parallelOut_955(v2c_out5[95]),
	.v2c_parallelOut_960(v2c_out0[96]),
	.v2c_parallelOut_961(v2c_out1[96]),
	.v2c_parallelOut_962(v2c_out2[96]),
	.v2c_parallelOut_963(v2c_out3[96]),
	.v2c_parallelOut_964(v2c_out4[96]),
	.v2c_parallelOut_965(v2c_out5[96]),
	.v2c_parallelOut_970(v2c_out0[97]),
	.v2c_parallelOut_971(v2c_out1[97]),
	.v2c_parallelOut_972(v2c_out2[97]),
	.v2c_parallelOut_973(v2c_out3[97]),
	.v2c_parallelOut_974(v2c_out4[97]),
	.v2c_parallelOut_975(v2c_out5[97]),
	.v2c_parallelOut_980(v2c_out0[98]),
	.v2c_parallelOut_981(v2c_out1[98]),
	.v2c_parallelOut_982(v2c_out2[98]),
	.v2c_parallelOut_983(v2c_out3[98]),
	.v2c_parallelOut_984(v2c_out4[98]),
	.v2c_parallelOut_985(v2c_out5[98]),
	.v2c_parallelOut_990(v2c_out0[99]),
	.v2c_parallelOut_991(v2c_out1[99]),
	.v2c_parallelOut_992(v2c_out2[99]),
	.v2c_parallelOut_993(v2c_out3[99]),
	.v2c_parallelOut_994(v2c_out4[99]),
	.v2c_parallelOut_995(v2c_out5[99]),
	.v2c_parallelOut_1000(v2c_out0[100]),
	.v2c_parallelOut_1001(v2c_out1[100]),
	.v2c_parallelOut_1002(v2c_out2[100]),
	.v2c_parallelOut_1003(v2c_out3[100]),
	.v2c_parallelOut_1004(v2c_out4[100]),
	.v2c_parallelOut_1005(v2c_out5[100]),
	.v2c_parallelOut_1010(v2c_out0[101]),
	.v2c_parallelOut_1011(v2c_out1[101]),
	.v2c_parallelOut_1012(v2c_out2[101]),
	.v2c_parallelOut_1013(v2c_out3[101]),
	.v2c_parallelOut_1014(v2c_out4[101]),
	.v2c_parallelOut_1015(v2c_out5[101]),
	
	// N number of check-to-Variable message buses, each of which is d_v bit width outgoing to serial-to-parallel converters
	.c2v_parallelOut_00(c2v_out0[0]),
	.c2v_parallelOut_01(c2v_out1[0]),
	.c2v_parallelOut_02(c2v_out2[0]),
	.c2v_parallelOut_10(c2v_out0[1]),
	.c2v_parallelOut_11(c2v_out1[1]),
	.c2v_parallelOut_12(c2v_out2[1]),
	.c2v_parallelOut_20(c2v_out0[2]),
	.c2v_parallelOut_21(c2v_out1[2]),
	.c2v_parallelOut_22(c2v_out2[2]),
	.c2v_parallelOut_30(c2v_out0[3]),
	.c2v_parallelOut_31(c2v_out1[3]),
	.c2v_parallelOut_32(c2v_out2[3]),
	.c2v_parallelOut_40(c2v_out0[4]),
	.c2v_parallelOut_41(c2v_out1[4]),
	.c2v_parallelOut_42(c2v_out2[4]),
	.c2v_parallelOut_50(c2v_out0[5]),
	.c2v_parallelOut_51(c2v_out1[5]),
	.c2v_parallelOut_52(c2v_out2[5]),
	.c2v_parallelOut_60(c2v_out0[6]),
	.c2v_parallelOut_61(c2v_out1[6]),
	.c2v_parallelOut_62(c2v_out2[6]),
	.c2v_parallelOut_70(c2v_out0[7]),
	.c2v_parallelOut_71(c2v_out1[7]),
	.c2v_parallelOut_72(c2v_out2[7]),
	.c2v_parallelOut_80(c2v_out0[8]),
	.c2v_parallelOut_81(c2v_out1[8]),
	.c2v_parallelOut_82(c2v_out2[8]),
	.c2v_parallelOut_90(c2v_out0[9]),
	.c2v_parallelOut_91(c2v_out1[9]),
	.c2v_parallelOut_92(c2v_out2[9]),
	.c2v_parallelOut_100(c2v_out0[10]),
	.c2v_parallelOut_101(c2v_out1[10]),
	.c2v_parallelOut_102(c2v_out2[10]),
	.c2v_parallelOut_110(c2v_out0[11]),
	.c2v_parallelOut_111(c2v_out1[11]),
	.c2v_parallelOut_112(c2v_out2[11]),
	.c2v_parallelOut_120(c2v_out0[12]),
	.c2v_parallelOut_121(c2v_out1[12]),
	.c2v_parallelOut_122(c2v_out2[12]),
	.c2v_parallelOut_130(c2v_out0[13]),
	.c2v_parallelOut_131(c2v_out1[13]),
	.c2v_parallelOut_132(c2v_out2[13]),
	.c2v_parallelOut_140(c2v_out0[14]),
	.c2v_parallelOut_141(c2v_out1[14]),
	.c2v_parallelOut_142(c2v_out2[14]),
	.c2v_parallelOut_150(c2v_out0[15]),
	.c2v_parallelOut_151(c2v_out1[15]),
	.c2v_parallelOut_152(c2v_out2[15]),
	.c2v_parallelOut_160(c2v_out0[16]),
	.c2v_parallelOut_161(c2v_out1[16]),
	.c2v_parallelOut_162(c2v_out2[16]),
	.c2v_parallelOut_170(c2v_out0[17]),
	.c2v_parallelOut_171(c2v_out1[17]),
	.c2v_parallelOut_172(c2v_out2[17]),
	.c2v_parallelOut_180(c2v_out0[18]),
	.c2v_parallelOut_181(c2v_out1[18]),
	.c2v_parallelOut_182(c2v_out2[18]),
	.c2v_parallelOut_190(c2v_out0[19]),
	.c2v_parallelOut_191(c2v_out1[19]),
	.c2v_parallelOut_192(c2v_out2[19]),
	.c2v_parallelOut_200(c2v_out0[20]),
	.c2v_parallelOut_201(c2v_out1[20]),
	.c2v_parallelOut_202(c2v_out2[20]),
	.c2v_parallelOut_210(c2v_out0[21]),
	.c2v_parallelOut_211(c2v_out1[21]),
	.c2v_parallelOut_212(c2v_out2[21]),
	.c2v_parallelOut_220(c2v_out0[22]),
	.c2v_parallelOut_221(c2v_out1[22]),
	.c2v_parallelOut_222(c2v_out2[22]),
	.c2v_parallelOut_230(c2v_out0[23]),
	.c2v_parallelOut_231(c2v_out1[23]),
	.c2v_parallelOut_232(c2v_out2[23]),
	.c2v_parallelOut_240(c2v_out0[24]),
	.c2v_parallelOut_241(c2v_out1[24]),
	.c2v_parallelOut_242(c2v_out2[24]),
	.c2v_parallelOut_250(c2v_out0[25]),
	.c2v_parallelOut_251(c2v_out1[25]),
	.c2v_parallelOut_252(c2v_out2[25]),
	.c2v_parallelOut_260(c2v_out0[26]),
	.c2v_parallelOut_261(c2v_out1[26]),
	.c2v_parallelOut_262(c2v_out2[26]),
	.c2v_parallelOut_270(c2v_out0[27]),
	.c2v_parallelOut_271(c2v_out1[27]),
	.c2v_parallelOut_272(c2v_out2[27]),
	.c2v_parallelOut_280(c2v_out0[28]),
	.c2v_parallelOut_281(c2v_out1[28]),
	.c2v_parallelOut_282(c2v_out2[28]),
	.c2v_parallelOut_290(c2v_out0[29]),
	.c2v_parallelOut_291(c2v_out1[29]),
	.c2v_parallelOut_292(c2v_out2[29]),
	.c2v_parallelOut_300(c2v_out0[30]),
	.c2v_parallelOut_301(c2v_out1[30]),
	.c2v_parallelOut_302(c2v_out2[30]),
	.c2v_parallelOut_310(c2v_out0[31]),
	.c2v_parallelOut_311(c2v_out1[31]),
	.c2v_parallelOut_312(c2v_out2[31]),
	.c2v_parallelOut_320(c2v_out0[32]),
	.c2v_parallelOut_321(c2v_out1[32]),
	.c2v_parallelOut_322(c2v_out2[32]),
	.c2v_parallelOut_330(c2v_out0[33]),
	.c2v_parallelOut_331(c2v_out1[33]),
	.c2v_parallelOut_332(c2v_out2[33]),
	.c2v_parallelOut_340(c2v_out0[34]),
	.c2v_parallelOut_341(c2v_out1[34]),
	.c2v_parallelOut_342(c2v_out2[34]),
	.c2v_parallelOut_350(c2v_out0[35]),
	.c2v_parallelOut_351(c2v_out1[35]),
	.c2v_parallelOut_352(c2v_out2[35]),
	.c2v_parallelOut_360(c2v_out0[36]),
	.c2v_parallelOut_361(c2v_out1[36]),
	.c2v_parallelOut_362(c2v_out2[36]),
	.c2v_parallelOut_370(c2v_out0[37]),
	.c2v_parallelOut_371(c2v_out1[37]),
	.c2v_parallelOut_372(c2v_out2[37]),
	.c2v_parallelOut_380(c2v_out0[38]),
	.c2v_parallelOut_381(c2v_out1[38]),
	.c2v_parallelOut_382(c2v_out2[38]),
	.c2v_parallelOut_390(c2v_out0[39]),
	.c2v_parallelOut_391(c2v_out1[39]),
	.c2v_parallelOut_392(c2v_out2[39]),
	.c2v_parallelOut_400(c2v_out0[40]),
	.c2v_parallelOut_401(c2v_out1[40]),
	.c2v_parallelOut_402(c2v_out2[40]),
	.c2v_parallelOut_410(c2v_out0[41]),
	.c2v_parallelOut_411(c2v_out1[41]),
	.c2v_parallelOut_412(c2v_out2[41]),
	.c2v_parallelOut_420(c2v_out0[42]),
	.c2v_parallelOut_421(c2v_out1[42]),
	.c2v_parallelOut_422(c2v_out2[42]),
	.c2v_parallelOut_430(c2v_out0[43]),
	.c2v_parallelOut_431(c2v_out1[43]),
	.c2v_parallelOut_432(c2v_out2[43]),
	.c2v_parallelOut_440(c2v_out0[44]),
	.c2v_parallelOut_441(c2v_out1[44]),
	.c2v_parallelOut_442(c2v_out2[44]),
	.c2v_parallelOut_450(c2v_out0[45]),
	.c2v_parallelOut_451(c2v_out1[45]),
	.c2v_parallelOut_452(c2v_out2[45]),
	.c2v_parallelOut_460(c2v_out0[46]),
	.c2v_parallelOut_461(c2v_out1[46]),
	.c2v_parallelOut_462(c2v_out2[46]),
	.c2v_parallelOut_470(c2v_out0[47]),
	.c2v_parallelOut_471(c2v_out1[47]),
	.c2v_parallelOut_472(c2v_out2[47]),
	.c2v_parallelOut_480(c2v_out0[48]),
	.c2v_parallelOut_481(c2v_out1[48]),
	.c2v_parallelOut_482(c2v_out2[48]),
	.c2v_parallelOut_490(c2v_out0[49]),
	.c2v_parallelOut_491(c2v_out1[49]),
	.c2v_parallelOut_492(c2v_out2[49]),
	.c2v_parallelOut_500(c2v_out0[50]),
	.c2v_parallelOut_501(c2v_out1[50]),
	.c2v_parallelOut_502(c2v_out2[50]),
	.c2v_parallelOut_510(c2v_out0[51]),
	.c2v_parallelOut_511(c2v_out1[51]),
	.c2v_parallelOut_512(c2v_out2[51]),
	.c2v_parallelOut_520(c2v_out0[52]),
	.c2v_parallelOut_521(c2v_out1[52]),
	.c2v_parallelOut_522(c2v_out2[52]),
	.c2v_parallelOut_530(c2v_out0[53]),
	.c2v_parallelOut_531(c2v_out1[53]),
	.c2v_parallelOut_532(c2v_out2[53]),
	.c2v_parallelOut_540(c2v_out0[54]),
	.c2v_parallelOut_541(c2v_out1[54]),
	.c2v_parallelOut_542(c2v_out2[54]),
	.c2v_parallelOut_550(c2v_out0[55]),
	.c2v_parallelOut_551(c2v_out1[55]),
	.c2v_parallelOut_552(c2v_out2[55]),
	.c2v_parallelOut_560(c2v_out0[56]),
	.c2v_parallelOut_561(c2v_out1[56]),
	.c2v_parallelOut_562(c2v_out2[56]),
	.c2v_parallelOut_570(c2v_out0[57]),
	.c2v_parallelOut_571(c2v_out1[57]),
	.c2v_parallelOut_572(c2v_out2[57]),
	.c2v_parallelOut_580(c2v_out0[58]),
	.c2v_parallelOut_581(c2v_out1[58]),
	.c2v_parallelOut_582(c2v_out2[58]),
	.c2v_parallelOut_590(c2v_out0[59]),
	.c2v_parallelOut_591(c2v_out1[59]),
	.c2v_parallelOut_592(c2v_out2[59]),
	.c2v_parallelOut_600(c2v_out0[60]),
	.c2v_parallelOut_601(c2v_out1[60]),
	.c2v_parallelOut_602(c2v_out2[60]),
	.c2v_parallelOut_610(c2v_out0[61]),
	.c2v_parallelOut_611(c2v_out1[61]),
	.c2v_parallelOut_612(c2v_out2[61]),
	.c2v_parallelOut_620(c2v_out0[62]),
	.c2v_parallelOut_621(c2v_out1[62]),
	.c2v_parallelOut_622(c2v_out2[62]),
	.c2v_parallelOut_630(c2v_out0[63]),
	.c2v_parallelOut_631(c2v_out1[63]),
	.c2v_parallelOut_632(c2v_out2[63]),
	.c2v_parallelOut_640(c2v_out0[64]),
	.c2v_parallelOut_641(c2v_out1[64]),
	.c2v_parallelOut_642(c2v_out2[64]),
	.c2v_parallelOut_650(c2v_out0[65]),
	.c2v_parallelOut_651(c2v_out1[65]),
	.c2v_parallelOut_652(c2v_out2[65]),
	.c2v_parallelOut_660(c2v_out0[66]),
	.c2v_parallelOut_661(c2v_out1[66]),
	.c2v_parallelOut_662(c2v_out2[66]),
	.c2v_parallelOut_670(c2v_out0[67]),
	.c2v_parallelOut_671(c2v_out1[67]),
	.c2v_parallelOut_672(c2v_out2[67]),
	.c2v_parallelOut_680(c2v_out0[68]),
	.c2v_parallelOut_681(c2v_out1[68]),
	.c2v_parallelOut_682(c2v_out2[68]),
	.c2v_parallelOut_690(c2v_out0[69]),
	.c2v_parallelOut_691(c2v_out1[69]),
	.c2v_parallelOut_692(c2v_out2[69]),
	.c2v_parallelOut_700(c2v_out0[70]),
	.c2v_parallelOut_701(c2v_out1[70]),
	.c2v_parallelOut_702(c2v_out2[70]),
	.c2v_parallelOut_710(c2v_out0[71]),
	.c2v_parallelOut_711(c2v_out1[71]),
	.c2v_parallelOut_712(c2v_out2[71]),
	.c2v_parallelOut_720(c2v_out0[72]),
	.c2v_parallelOut_721(c2v_out1[72]),
	.c2v_parallelOut_722(c2v_out2[72]),
	.c2v_parallelOut_730(c2v_out0[73]),
	.c2v_parallelOut_731(c2v_out1[73]),
	.c2v_parallelOut_732(c2v_out2[73]),
	.c2v_parallelOut_740(c2v_out0[74]),
	.c2v_parallelOut_741(c2v_out1[74]),
	.c2v_parallelOut_742(c2v_out2[74]),
	.c2v_parallelOut_750(c2v_out0[75]),
	.c2v_parallelOut_751(c2v_out1[75]),
	.c2v_parallelOut_752(c2v_out2[75]),
	.c2v_parallelOut_760(c2v_out0[76]),
	.c2v_parallelOut_761(c2v_out1[76]),
	.c2v_parallelOut_762(c2v_out2[76]),
	.c2v_parallelOut_770(c2v_out0[77]),
	.c2v_parallelOut_771(c2v_out1[77]),
	.c2v_parallelOut_772(c2v_out2[77]),
	.c2v_parallelOut_780(c2v_out0[78]),
	.c2v_parallelOut_781(c2v_out1[78]),
	.c2v_parallelOut_782(c2v_out2[78]),
	.c2v_parallelOut_790(c2v_out0[79]),
	.c2v_parallelOut_791(c2v_out1[79]),
	.c2v_parallelOut_792(c2v_out2[79]),
	.c2v_parallelOut_800(c2v_out0[80]),
	.c2v_parallelOut_801(c2v_out1[80]),
	.c2v_parallelOut_802(c2v_out2[80]),
	.c2v_parallelOut_810(c2v_out0[81]),
	.c2v_parallelOut_811(c2v_out1[81]),
	.c2v_parallelOut_812(c2v_out2[81]),
	.c2v_parallelOut_820(c2v_out0[82]),
	.c2v_parallelOut_821(c2v_out1[82]),
	.c2v_parallelOut_822(c2v_out2[82]),
	.c2v_parallelOut_830(c2v_out0[83]),
	.c2v_parallelOut_831(c2v_out1[83]),
	.c2v_parallelOut_832(c2v_out2[83]),
	.c2v_parallelOut_840(c2v_out0[84]),
	.c2v_parallelOut_841(c2v_out1[84]),
	.c2v_parallelOut_842(c2v_out2[84]),
	.c2v_parallelOut_850(c2v_out0[85]),
	.c2v_parallelOut_851(c2v_out1[85]),
	.c2v_parallelOut_852(c2v_out2[85]),
	.c2v_parallelOut_860(c2v_out0[86]),
	.c2v_parallelOut_861(c2v_out1[86]),
	.c2v_parallelOut_862(c2v_out2[86]),
	.c2v_parallelOut_870(c2v_out0[87]),
	.c2v_parallelOut_871(c2v_out1[87]),
	.c2v_parallelOut_872(c2v_out2[87]),
	.c2v_parallelOut_880(c2v_out0[88]),
	.c2v_parallelOut_881(c2v_out1[88]),
	.c2v_parallelOut_882(c2v_out2[88]),
	.c2v_parallelOut_890(c2v_out0[89]),
	.c2v_parallelOut_891(c2v_out1[89]),
	.c2v_parallelOut_892(c2v_out2[89]),
	.c2v_parallelOut_900(c2v_out0[90]),
	.c2v_parallelOut_901(c2v_out1[90]),
	.c2v_parallelOut_902(c2v_out2[90]),
	.c2v_parallelOut_910(c2v_out0[91]),
	.c2v_parallelOut_911(c2v_out1[91]),
	.c2v_parallelOut_912(c2v_out2[91]),
	.c2v_parallelOut_920(c2v_out0[92]),
	.c2v_parallelOut_921(c2v_out1[92]),
	.c2v_parallelOut_922(c2v_out2[92]),
	.c2v_parallelOut_930(c2v_out0[93]),
	.c2v_parallelOut_931(c2v_out1[93]),
	.c2v_parallelOut_932(c2v_out2[93]),
	.c2v_parallelOut_940(c2v_out0[94]),
	.c2v_parallelOut_941(c2v_out1[94]),
	.c2v_parallelOut_942(c2v_out2[94]),
	.c2v_parallelOut_950(c2v_out0[95]),
	.c2v_parallelOut_951(c2v_out1[95]),
	.c2v_parallelOut_952(c2v_out2[95]),
	.c2v_parallelOut_960(c2v_out0[96]),
	.c2v_parallelOut_961(c2v_out1[96]),
	.c2v_parallelOut_962(c2v_out2[96]),
	.c2v_parallelOut_970(c2v_out0[97]),
	.c2v_parallelOut_971(c2v_out1[97]),
	.c2v_parallelOut_972(c2v_out2[97]),
	.c2v_parallelOut_980(c2v_out0[98]),
	.c2v_parallelOut_981(c2v_out1[98]),
	.c2v_parallelOut_982(c2v_out2[98]),
	.c2v_parallelOut_990(c2v_out0[99]),
	.c2v_parallelOut_991(c2v_out1[99]),
	.c2v_parallelOut_992(c2v_out2[99]),
	.c2v_parallelOut_1000(c2v_out0[100]),
	.c2v_parallelOut_1001(c2v_out1[100]),
	.c2v_parallelOut_1002(c2v_out2[100]),
	.c2v_parallelOut_1010(c2v_out0[101]),
	.c2v_parallelOut_1011(c2v_out1[101]),
	.c2v_parallelOut_1012(c2v_out2[101]),
	.c2v_parallelOut_1020(c2v_out0[102]),
	.c2v_parallelOut_1021(c2v_out1[102]),
	.c2v_parallelOut_1022(c2v_out2[102]),
	.c2v_parallelOut_1030(c2v_out0[103]),
	.c2v_parallelOut_1031(c2v_out1[103]),
	.c2v_parallelOut_1032(c2v_out2[103]),
	.c2v_parallelOut_1040(c2v_out0[104]),
	.c2v_parallelOut_1041(c2v_out1[104]),
	.c2v_parallelOut_1042(c2v_out2[104]),
	.c2v_parallelOut_1050(c2v_out0[105]),
	.c2v_parallelOut_1051(c2v_out1[105]),
	.c2v_parallelOut_1052(c2v_out2[105]),
	.c2v_parallelOut_1060(c2v_out0[106]),
	.c2v_parallelOut_1061(c2v_out1[106]),
	.c2v_parallelOut_1062(c2v_out2[106]),
	.c2v_parallelOut_1070(c2v_out0[107]),
	.c2v_parallelOut_1071(c2v_out1[107]),
	.c2v_parallelOut_1072(c2v_out2[107]),
	.c2v_parallelOut_1080(c2v_out0[108]),
	.c2v_parallelOut_1081(c2v_out1[108]),
	.c2v_parallelOut_1082(c2v_out2[108]),
	.c2v_parallelOut_1090(c2v_out0[109]),
	.c2v_parallelOut_1091(c2v_out1[109]),
	.c2v_parallelOut_1092(c2v_out2[109]),
	.c2v_parallelOut_1100(c2v_out0[110]),
	.c2v_parallelOut_1101(c2v_out1[110]),
	.c2v_parallelOut_1102(c2v_out2[110]),
	.c2v_parallelOut_1110(c2v_out0[111]),
	.c2v_parallelOut_1111(c2v_out1[111]),
	.c2v_parallelOut_1112(c2v_out2[111]),
	.c2v_parallelOut_1120(c2v_out0[112]),
	.c2v_parallelOut_1121(c2v_out1[112]),
	.c2v_parallelOut_1122(c2v_out2[112]),
	.c2v_parallelOut_1130(c2v_out0[113]),
	.c2v_parallelOut_1131(c2v_out1[113]),
	.c2v_parallelOut_1132(c2v_out2[113]),
	.c2v_parallelOut_1140(c2v_out0[114]),
	.c2v_parallelOut_1141(c2v_out1[114]),
	.c2v_parallelOut_1142(c2v_out2[114]),
	.c2v_parallelOut_1150(c2v_out0[115]),
	.c2v_parallelOut_1151(c2v_out1[115]),
	.c2v_parallelOut_1152(c2v_out2[115]),
	.c2v_parallelOut_1160(c2v_out0[116]),
	.c2v_parallelOut_1161(c2v_out1[116]),
	.c2v_parallelOut_1162(c2v_out2[116]),
	.c2v_parallelOut_1170(c2v_out0[117]),
	.c2v_parallelOut_1171(c2v_out1[117]),
	.c2v_parallelOut_1172(c2v_out2[117]),
	.c2v_parallelOut_1180(c2v_out0[118]),
	.c2v_parallelOut_1181(c2v_out1[118]),
	.c2v_parallelOut_1182(c2v_out2[118]),
	.c2v_parallelOut_1190(c2v_out0[119]),
	.c2v_parallelOut_1191(c2v_out1[119]),
	.c2v_parallelOut_1192(c2v_out2[119]),
	.c2v_parallelOut_1200(c2v_out0[120]),
	.c2v_parallelOut_1201(c2v_out1[120]),
	.c2v_parallelOut_1202(c2v_out2[120]),
	.c2v_parallelOut_1210(c2v_out0[121]),
	.c2v_parallelOut_1211(c2v_out1[121]),
	.c2v_parallelOut_1212(c2v_out2[121]),
	.c2v_parallelOut_1220(c2v_out0[122]),
	.c2v_parallelOut_1221(c2v_out1[122]),
	.c2v_parallelOut_1222(c2v_out2[122]),
	.c2v_parallelOut_1230(c2v_out0[123]),
	.c2v_parallelOut_1231(c2v_out1[123]),
	.c2v_parallelOut_1232(c2v_out2[123]),
	.c2v_parallelOut_1240(c2v_out0[124]),
	.c2v_parallelOut_1241(c2v_out1[124]),
	.c2v_parallelOut_1242(c2v_out2[124]),
	.c2v_parallelOut_1250(c2v_out0[125]),
	.c2v_parallelOut_1251(c2v_out1[125]),
	.c2v_parallelOut_1252(c2v_out2[125]),
	.c2v_parallelOut_1260(c2v_out0[126]),
	.c2v_parallelOut_1261(c2v_out1[126]),
	.c2v_parallelOut_1262(c2v_out2[126]),
	.c2v_parallelOut_1270(c2v_out0[127]),
	.c2v_parallelOut_1271(c2v_out1[127]),
	.c2v_parallelOut_1272(c2v_out2[127]),
	.c2v_parallelOut_1280(c2v_out0[128]),
	.c2v_parallelOut_1281(c2v_out1[128]),
	.c2v_parallelOut_1282(c2v_out2[128]),
	.c2v_parallelOut_1290(c2v_out0[129]),
	.c2v_parallelOut_1291(c2v_out1[129]),
	.c2v_parallelOut_1292(c2v_out2[129]),
	.c2v_parallelOut_1300(c2v_out0[130]),
	.c2v_parallelOut_1301(c2v_out1[130]),
	.c2v_parallelOut_1302(c2v_out2[130]),
	.c2v_parallelOut_1310(c2v_out0[131]),
	.c2v_parallelOut_1311(c2v_out1[131]),
	.c2v_parallelOut_1312(c2v_out2[131]),
	.c2v_parallelOut_1320(c2v_out0[132]),
	.c2v_parallelOut_1321(c2v_out1[132]),
	.c2v_parallelOut_1322(c2v_out2[132]),
	.c2v_parallelOut_1330(c2v_out0[133]),
	.c2v_parallelOut_1331(c2v_out1[133]),
	.c2v_parallelOut_1332(c2v_out2[133]),
	.c2v_parallelOut_1340(c2v_out0[134]),
	.c2v_parallelOut_1341(c2v_out1[134]),
	.c2v_parallelOut_1342(c2v_out2[134]),
	.c2v_parallelOut_1350(c2v_out0[135]),
	.c2v_parallelOut_1351(c2v_out1[135]),
	.c2v_parallelOut_1352(c2v_out2[135]),
	.c2v_parallelOut_1360(c2v_out0[136]),
	.c2v_parallelOut_1361(c2v_out1[136]),
	.c2v_parallelOut_1362(c2v_out2[136]),
	.c2v_parallelOut_1370(c2v_out0[137]),
	.c2v_parallelOut_1371(c2v_out1[137]),
	.c2v_parallelOut_1372(c2v_out2[137]),
	.c2v_parallelOut_1380(c2v_out0[138]),
	.c2v_parallelOut_1381(c2v_out1[138]),
	.c2v_parallelOut_1382(c2v_out2[138]),
	.c2v_parallelOut_1390(c2v_out0[139]),
	.c2v_parallelOut_1391(c2v_out1[139]),
	.c2v_parallelOut_1392(c2v_out2[139]),
	.c2v_parallelOut_1400(c2v_out0[140]),
	.c2v_parallelOut_1401(c2v_out1[140]),
	.c2v_parallelOut_1402(c2v_out2[140]),
	.c2v_parallelOut_1410(c2v_out0[141]),
	.c2v_parallelOut_1411(c2v_out1[141]),
	.c2v_parallelOut_1412(c2v_out2[141]),
	.c2v_parallelOut_1420(c2v_out0[142]),
	.c2v_parallelOut_1421(c2v_out1[142]),
	.c2v_parallelOut_1422(c2v_out2[142]),
	.c2v_parallelOut_1430(c2v_out0[143]),
	.c2v_parallelOut_1431(c2v_out1[143]),
	.c2v_parallelOut_1432(c2v_out2[143]),
	.c2v_parallelOut_1440(c2v_out0[144]),
	.c2v_parallelOut_1441(c2v_out1[144]),
	.c2v_parallelOut_1442(c2v_out2[144]),
	.c2v_parallelOut_1450(c2v_out0[145]),
	.c2v_parallelOut_1451(c2v_out1[145]),
	.c2v_parallelOut_1452(c2v_out2[145]),
	.c2v_parallelOut_1460(c2v_out0[146]),
	.c2v_parallelOut_1461(c2v_out1[146]),
	.c2v_parallelOut_1462(c2v_out2[146]),
	.c2v_parallelOut_1470(c2v_out0[147]),
	.c2v_parallelOut_1471(c2v_out1[147]),
	.c2v_parallelOut_1472(c2v_out2[147]),
	.c2v_parallelOut_1480(c2v_out0[148]),
	.c2v_parallelOut_1481(c2v_out1[148]),
	.c2v_parallelOut_1482(c2v_out2[148]),
	.c2v_parallelOut_1490(c2v_out0[149]),
	.c2v_parallelOut_1491(c2v_out1[149]),
	.c2v_parallelOut_1492(c2v_out2[149]),
	.c2v_parallelOut_1500(c2v_out0[150]),
	.c2v_parallelOut_1501(c2v_out1[150]),
	.c2v_parallelOut_1502(c2v_out2[150]),
	.c2v_parallelOut_1510(c2v_out0[151]),
	.c2v_parallelOut_1511(c2v_out1[151]),
	.c2v_parallelOut_1512(c2v_out2[151]),
	.c2v_parallelOut_1520(c2v_out0[152]),
	.c2v_parallelOut_1521(c2v_out1[152]),
	.c2v_parallelOut_1522(c2v_out2[152]),
	.c2v_parallelOut_1530(c2v_out0[153]),
	.c2v_parallelOut_1531(c2v_out1[153]),
	.c2v_parallelOut_1532(c2v_out2[153]),
	.c2v_parallelOut_1540(c2v_out0[154]),
	.c2v_parallelOut_1541(c2v_out1[154]),
	.c2v_parallelOut_1542(c2v_out2[154]),
	.c2v_parallelOut_1550(c2v_out0[155]),
	.c2v_parallelOut_1551(c2v_out1[155]),
	.c2v_parallelOut_1552(c2v_out2[155]),
	.c2v_parallelOut_1560(c2v_out0[156]),
	.c2v_parallelOut_1561(c2v_out1[156]),
	.c2v_parallelOut_1562(c2v_out2[156]),
	.c2v_parallelOut_1570(c2v_out0[157]),
	.c2v_parallelOut_1571(c2v_out1[157]),
	.c2v_parallelOut_1572(c2v_out2[157]),
	.c2v_parallelOut_1580(c2v_out0[158]),
	.c2v_parallelOut_1581(c2v_out1[158]),
	.c2v_parallelOut_1582(c2v_out2[158]),
	.c2v_parallelOut_1590(c2v_out0[159]),
	.c2v_parallelOut_1591(c2v_out1[159]),
	.c2v_parallelOut_1592(c2v_out2[159]),
	.c2v_parallelOut_1600(c2v_out0[160]),
	.c2v_parallelOut_1601(c2v_out1[160]),
	.c2v_parallelOut_1602(c2v_out2[160]),
	.c2v_parallelOut_1610(c2v_out0[161]),
	.c2v_parallelOut_1611(c2v_out1[161]),
	.c2v_parallelOut_1612(c2v_out2[161]),
	.c2v_parallelOut_1620(c2v_out0[162]),
	.c2v_parallelOut_1621(c2v_out1[162]),
	.c2v_parallelOut_1622(c2v_out2[162]),
	.c2v_parallelOut_1630(c2v_out0[163]),
	.c2v_parallelOut_1631(c2v_out1[163]),
	.c2v_parallelOut_1632(c2v_out2[163]),
	.c2v_parallelOut_1640(c2v_out0[164]),
	.c2v_parallelOut_1641(c2v_out1[164]),
	.c2v_parallelOut_1642(c2v_out2[164]),
	.c2v_parallelOut_1650(c2v_out0[165]),
	.c2v_parallelOut_1651(c2v_out1[165]),
	.c2v_parallelOut_1652(c2v_out2[165]),
	.c2v_parallelOut_1660(c2v_out0[166]),
	.c2v_parallelOut_1661(c2v_out1[166]),
	.c2v_parallelOut_1662(c2v_out2[166]),
	.c2v_parallelOut_1670(c2v_out0[167]),
	.c2v_parallelOut_1671(c2v_out1[167]),
	.c2v_parallelOut_1672(c2v_out2[167]),
	.c2v_parallelOut_1680(c2v_out0[168]),
	.c2v_parallelOut_1681(c2v_out1[168]),
	.c2v_parallelOut_1682(c2v_out2[168]),
	.c2v_parallelOut_1690(c2v_out0[169]),
	.c2v_parallelOut_1691(c2v_out1[169]),
	.c2v_parallelOut_1692(c2v_out2[169]),
	.c2v_parallelOut_1700(c2v_out0[170]),
	.c2v_parallelOut_1701(c2v_out1[170]),
	.c2v_parallelOut_1702(c2v_out2[170]),
	.c2v_parallelOut_1710(c2v_out0[171]),
	.c2v_parallelOut_1711(c2v_out1[171]),
	.c2v_parallelOut_1712(c2v_out2[171]),
	.c2v_parallelOut_1720(c2v_out0[172]),
	.c2v_parallelOut_1721(c2v_out1[172]),
	.c2v_parallelOut_1722(c2v_out2[172]),
	.c2v_parallelOut_1730(c2v_out0[173]),
	.c2v_parallelOut_1731(c2v_out1[173]),
	.c2v_parallelOut_1732(c2v_out2[173]),
	.c2v_parallelOut_1740(c2v_out0[174]),
	.c2v_parallelOut_1741(c2v_out1[174]),
	.c2v_parallelOut_1742(c2v_out2[174]),
	.c2v_parallelOut_1750(c2v_out0[175]),
	.c2v_parallelOut_1751(c2v_out1[175]),
	.c2v_parallelOut_1752(c2v_out2[175]),
	.c2v_parallelOut_1760(c2v_out0[176]),
	.c2v_parallelOut_1761(c2v_out1[176]),
	.c2v_parallelOut_1762(c2v_out2[176]),
	.c2v_parallelOut_1770(c2v_out0[177]),
	.c2v_parallelOut_1771(c2v_out1[177]),
	.c2v_parallelOut_1772(c2v_out2[177]),
	.c2v_parallelOut_1780(c2v_out0[178]),
	.c2v_parallelOut_1781(c2v_out1[178]),
	.c2v_parallelOut_1782(c2v_out2[178]),
	.c2v_parallelOut_1790(c2v_out0[179]),
	.c2v_parallelOut_1791(c2v_out1[179]),
	.c2v_parallelOut_1792(c2v_out2[179]),
	.c2v_parallelOut_1800(c2v_out0[180]),
	.c2v_parallelOut_1801(c2v_out1[180]),
	.c2v_parallelOut_1802(c2v_out2[180]),
	.c2v_parallelOut_1810(c2v_out0[181]),
	.c2v_parallelOut_1811(c2v_out1[181]),
	.c2v_parallelOut_1812(c2v_out2[181]),
	.c2v_parallelOut_1820(c2v_out0[182]),
	.c2v_parallelOut_1821(c2v_out1[182]),
	.c2v_parallelOut_1822(c2v_out2[182]),
	.c2v_parallelOut_1830(c2v_out0[183]),
	.c2v_parallelOut_1831(c2v_out1[183]),
	.c2v_parallelOut_1832(c2v_out2[183]),
	.c2v_parallelOut_1840(c2v_out0[184]),
	.c2v_parallelOut_1841(c2v_out1[184]),
	.c2v_parallelOut_1842(c2v_out2[184]),
	.c2v_parallelOut_1850(c2v_out0[185]),
	.c2v_parallelOut_1851(c2v_out1[185]),
	.c2v_parallelOut_1852(c2v_out2[185]),
	.c2v_parallelOut_1860(c2v_out0[186]),
	.c2v_parallelOut_1861(c2v_out1[186]),
	.c2v_parallelOut_1862(c2v_out2[186]),
	.c2v_parallelOut_1870(c2v_out0[187]),
	.c2v_parallelOut_1871(c2v_out1[187]),
	.c2v_parallelOut_1872(c2v_out2[187]),
	.c2v_parallelOut_1880(c2v_out0[188]),
	.c2v_parallelOut_1881(c2v_out1[188]),
	.c2v_parallelOut_1882(c2v_out2[188]),
	.c2v_parallelOut_1890(c2v_out0[189]),
	.c2v_parallelOut_1891(c2v_out1[189]),
	.c2v_parallelOut_1892(c2v_out2[189]),
	.c2v_parallelOut_1900(c2v_out0[190]),
	.c2v_parallelOut_1901(c2v_out1[190]),
	.c2v_parallelOut_1902(c2v_out2[190]),
	.c2v_parallelOut_1910(c2v_out0[191]),
	.c2v_parallelOut_1911(c2v_out1[191]),
	.c2v_parallelOut_1912(c2v_out2[191]),
	.c2v_parallelOut_1920(c2v_out0[192]),
	.c2v_parallelOut_1921(c2v_out1[192]),
	.c2v_parallelOut_1922(c2v_out2[192]),
	.c2v_parallelOut_1930(c2v_out0[193]),
	.c2v_parallelOut_1931(c2v_out1[193]),
	.c2v_parallelOut_1932(c2v_out2[193]),
	.c2v_parallelOut_1940(c2v_out0[194]),
	.c2v_parallelOut_1941(c2v_out1[194]),
	.c2v_parallelOut_1942(c2v_out2[194]),
	.c2v_parallelOut_1950(c2v_out0[195]),
	.c2v_parallelOut_1951(c2v_out1[195]),
	.c2v_parallelOut_1952(c2v_out2[195]),
	.c2v_parallelOut_1960(c2v_out0[196]),
	.c2v_parallelOut_1961(c2v_out1[196]),
	.c2v_parallelOut_1962(c2v_out2[196]),
	.c2v_parallelOut_1970(c2v_out0[197]),
	.c2v_parallelOut_1971(c2v_out1[197]),
	.c2v_parallelOut_1972(c2v_out2[197]),
	.c2v_parallelOut_1980(c2v_out0[198]),
	.c2v_parallelOut_1981(c2v_out1[198]),
	.c2v_parallelOut_1982(c2v_out2[198]),
	.c2v_parallelOut_1990(c2v_out0[199]),
	.c2v_parallelOut_1991(c2v_out1[199]),
	.c2v_parallelOut_1992(c2v_out2[199]),
	.c2v_parallelOut_2000(c2v_out0[200]),
	.c2v_parallelOut_2001(c2v_out1[200]),
	.c2v_parallelOut_2002(c2v_out2[200]),
	.c2v_parallelOut_2010(c2v_out0[201]),
	.c2v_parallelOut_2011(c2v_out1[201]),
	.c2v_parallelOut_2012(c2v_out2[201]),
	.c2v_parallelOut_2020(c2v_out0[202]),
	.c2v_parallelOut_2021(c2v_out1[202]),
	.c2v_parallelOut_2022(c2v_out2[202]),
	.c2v_parallelOut_2030(c2v_out0[203]),
	.c2v_parallelOut_2031(c2v_out1[203]),
	.c2v_parallelOut_2032(c2v_out2[203]),
	
	.c2v_parallelIn_00(c2v_in0[0]),
	.c2v_parallelIn_01(c2v_in1[0]),
	.c2v_parallelIn_02(c2v_in2[0]),
	.c2v_parallelIn_03(c2v_in3[0]),
	.c2v_parallelIn_04(c2v_in4[0]),
	.c2v_parallelIn_05(c2v_in5[0]),
	.c2v_parallelIn_10(c2v_in0[1]),
	.c2v_parallelIn_11(c2v_in1[1]),
	.c2v_parallelIn_12(c2v_in2[1]),
	.c2v_parallelIn_13(c2v_in3[1]),
	.c2v_parallelIn_14(c2v_in4[1]),
	.c2v_parallelIn_15(c2v_in5[1]),
	.c2v_parallelIn_20(c2v_in0[2]),
	.c2v_parallelIn_21(c2v_in1[2]),
	.c2v_parallelIn_22(c2v_in2[2]),
	.c2v_parallelIn_23(c2v_in3[2]),
	.c2v_parallelIn_24(c2v_in4[2]),
	.c2v_parallelIn_25(c2v_in5[2]),
	.c2v_parallelIn_30(c2v_in0[3]),
	.c2v_parallelIn_31(c2v_in1[3]),
	.c2v_parallelIn_32(c2v_in2[3]),
	.c2v_parallelIn_33(c2v_in3[3]),
	.c2v_parallelIn_34(c2v_in4[3]),
	.c2v_parallelIn_35(c2v_in5[3]),
	.c2v_parallelIn_40(c2v_in0[4]),
	.c2v_parallelIn_41(c2v_in1[4]),
	.c2v_parallelIn_42(c2v_in2[4]),
	.c2v_parallelIn_43(c2v_in3[4]),
	.c2v_parallelIn_44(c2v_in4[4]),
	.c2v_parallelIn_45(c2v_in5[4]),
	.c2v_parallelIn_50(c2v_in0[5]),
	.c2v_parallelIn_51(c2v_in1[5]),
	.c2v_parallelIn_52(c2v_in2[5]),
	.c2v_parallelIn_53(c2v_in3[5]),
	.c2v_parallelIn_54(c2v_in4[5]),
	.c2v_parallelIn_55(c2v_in5[5]),
	.c2v_parallelIn_60(c2v_in0[6]),
	.c2v_parallelIn_61(c2v_in1[6]),
	.c2v_parallelIn_62(c2v_in2[6]),
	.c2v_parallelIn_63(c2v_in3[6]),
	.c2v_parallelIn_64(c2v_in4[6]),
	.c2v_parallelIn_65(c2v_in5[6]),
	.c2v_parallelIn_70(c2v_in0[7]),
	.c2v_parallelIn_71(c2v_in1[7]),
	.c2v_parallelIn_72(c2v_in2[7]),
	.c2v_parallelIn_73(c2v_in3[7]),
	.c2v_parallelIn_74(c2v_in4[7]),
	.c2v_parallelIn_75(c2v_in5[7]),
	.c2v_parallelIn_80(c2v_in0[8]),
	.c2v_parallelIn_81(c2v_in1[8]),
	.c2v_parallelIn_82(c2v_in2[8]),
	.c2v_parallelIn_83(c2v_in3[8]),
	.c2v_parallelIn_84(c2v_in4[8]),
	.c2v_parallelIn_85(c2v_in5[8]),
	.c2v_parallelIn_90(c2v_in0[9]),
	.c2v_parallelIn_91(c2v_in1[9]),
	.c2v_parallelIn_92(c2v_in2[9]),
	.c2v_parallelIn_93(c2v_in3[9]),
	.c2v_parallelIn_94(c2v_in4[9]),
	.c2v_parallelIn_95(c2v_in5[9]),
	.c2v_parallelIn_100(c2v_in0[10]),
	.c2v_parallelIn_101(c2v_in1[10]),
	.c2v_parallelIn_102(c2v_in2[10]),
	.c2v_parallelIn_103(c2v_in3[10]),
	.c2v_parallelIn_104(c2v_in4[10]),
	.c2v_parallelIn_105(c2v_in5[10]),
	.c2v_parallelIn_110(c2v_in0[11]),
	.c2v_parallelIn_111(c2v_in1[11]),
	.c2v_parallelIn_112(c2v_in2[11]),
	.c2v_parallelIn_113(c2v_in3[11]),
	.c2v_parallelIn_114(c2v_in4[11]),
	.c2v_parallelIn_115(c2v_in5[11]),
	.c2v_parallelIn_120(c2v_in0[12]),
	.c2v_parallelIn_121(c2v_in1[12]),
	.c2v_parallelIn_122(c2v_in2[12]),
	.c2v_parallelIn_123(c2v_in3[12]),
	.c2v_parallelIn_124(c2v_in4[12]),
	.c2v_parallelIn_125(c2v_in5[12]),
	.c2v_parallelIn_130(c2v_in0[13]),
	.c2v_parallelIn_131(c2v_in1[13]),
	.c2v_parallelIn_132(c2v_in2[13]),
	.c2v_parallelIn_133(c2v_in3[13]),
	.c2v_parallelIn_134(c2v_in4[13]),
	.c2v_parallelIn_135(c2v_in5[13]),
	.c2v_parallelIn_140(c2v_in0[14]),
	.c2v_parallelIn_141(c2v_in1[14]),
	.c2v_parallelIn_142(c2v_in2[14]),
	.c2v_parallelIn_143(c2v_in3[14]),
	.c2v_parallelIn_144(c2v_in4[14]),
	.c2v_parallelIn_145(c2v_in5[14]),
	.c2v_parallelIn_150(c2v_in0[15]),
	.c2v_parallelIn_151(c2v_in1[15]),
	.c2v_parallelIn_152(c2v_in2[15]),
	.c2v_parallelIn_153(c2v_in3[15]),
	.c2v_parallelIn_154(c2v_in4[15]),
	.c2v_parallelIn_155(c2v_in5[15]),
	.c2v_parallelIn_160(c2v_in0[16]),
	.c2v_parallelIn_161(c2v_in1[16]),
	.c2v_parallelIn_162(c2v_in2[16]),
	.c2v_parallelIn_163(c2v_in3[16]),
	.c2v_parallelIn_164(c2v_in4[16]),
	.c2v_parallelIn_165(c2v_in5[16]),
	.c2v_parallelIn_170(c2v_in0[17]),
	.c2v_parallelIn_171(c2v_in1[17]),
	.c2v_parallelIn_172(c2v_in2[17]),
	.c2v_parallelIn_173(c2v_in3[17]),
	.c2v_parallelIn_174(c2v_in4[17]),
	.c2v_parallelIn_175(c2v_in5[17]),
	.c2v_parallelIn_180(c2v_in0[18]),
	.c2v_parallelIn_181(c2v_in1[18]),
	.c2v_parallelIn_182(c2v_in2[18]),
	.c2v_parallelIn_183(c2v_in3[18]),
	.c2v_parallelIn_184(c2v_in4[18]),
	.c2v_parallelIn_185(c2v_in5[18]),
	.c2v_parallelIn_190(c2v_in0[19]),
	.c2v_parallelIn_191(c2v_in1[19]),
	.c2v_parallelIn_192(c2v_in2[19]),
	.c2v_parallelIn_193(c2v_in3[19]),
	.c2v_parallelIn_194(c2v_in4[19]),
	.c2v_parallelIn_195(c2v_in5[19]),
	.c2v_parallelIn_200(c2v_in0[20]),
	.c2v_parallelIn_201(c2v_in1[20]),
	.c2v_parallelIn_202(c2v_in2[20]),
	.c2v_parallelIn_203(c2v_in3[20]),
	.c2v_parallelIn_204(c2v_in4[20]),
	.c2v_parallelIn_205(c2v_in5[20]),
	.c2v_parallelIn_210(c2v_in0[21]),
	.c2v_parallelIn_211(c2v_in1[21]),
	.c2v_parallelIn_212(c2v_in2[21]),
	.c2v_parallelIn_213(c2v_in3[21]),
	.c2v_parallelIn_214(c2v_in4[21]),
	.c2v_parallelIn_215(c2v_in5[21]),
	.c2v_parallelIn_220(c2v_in0[22]),
	.c2v_parallelIn_221(c2v_in1[22]),
	.c2v_parallelIn_222(c2v_in2[22]),
	.c2v_parallelIn_223(c2v_in3[22]),
	.c2v_parallelIn_224(c2v_in4[22]),
	.c2v_parallelIn_225(c2v_in5[22]),
	.c2v_parallelIn_230(c2v_in0[23]),
	.c2v_parallelIn_231(c2v_in1[23]),
	.c2v_parallelIn_232(c2v_in2[23]),
	.c2v_parallelIn_233(c2v_in3[23]),
	.c2v_parallelIn_234(c2v_in4[23]),
	.c2v_parallelIn_235(c2v_in5[23]),
	.c2v_parallelIn_240(c2v_in0[24]),
	.c2v_parallelIn_241(c2v_in1[24]),
	.c2v_parallelIn_242(c2v_in2[24]),
	.c2v_parallelIn_243(c2v_in3[24]),
	.c2v_parallelIn_244(c2v_in4[24]),
	.c2v_parallelIn_245(c2v_in5[24]),
	.c2v_parallelIn_250(c2v_in0[25]),
	.c2v_parallelIn_251(c2v_in1[25]),
	.c2v_parallelIn_252(c2v_in2[25]),
	.c2v_parallelIn_253(c2v_in3[25]),
	.c2v_parallelIn_254(c2v_in4[25]),
	.c2v_parallelIn_255(c2v_in5[25]),
	.c2v_parallelIn_260(c2v_in0[26]),
	.c2v_parallelIn_261(c2v_in1[26]),
	.c2v_parallelIn_262(c2v_in2[26]),
	.c2v_parallelIn_263(c2v_in3[26]),
	.c2v_parallelIn_264(c2v_in4[26]),
	.c2v_parallelIn_265(c2v_in5[26]),
	.c2v_parallelIn_270(c2v_in0[27]),
	.c2v_parallelIn_271(c2v_in1[27]),
	.c2v_parallelIn_272(c2v_in2[27]),
	.c2v_parallelIn_273(c2v_in3[27]),
	.c2v_parallelIn_274(c2v_in4[27]),
	.c2v_parallelIn_275(c2v_in5[27]),
	.c2v_parallelIn_280(c2v_in0[28]),
	.c2v_parallelIn_281(c2v_in1[28]),
	.c2v_parallelIn_282(c2v_in2[28]),
	.c2v_parallelIn_283(c2v_in3[28]),
	.c2v_parallelIn_284(c2v_in4[28]),
	.c2v_parallelIn_285(c2v_in5[28]),
	.c2v_parallelIn_290(c2v_in0[29]),
	.c2v_parallelIn_291(c2v_in1[29]),
	.c2v_parallelIn_292(c2v_in2[29]),
	.c2v_parallelIn_293(c2v_in3[29]),
	.c2v_parallelIn_294(c2v_in4[29]),
	.c2v_parallelIn_295(c2v_in5[29]),
	.c2v_parallelIn_300(c2v_in0[30]),
	.c2v_parallelIn_301(c2v_in1[30]),
	.c2v_parallelIn_302(c2v_in2[30]),
	.c2v_parallelIn_303(c2v_in3[30]),
	.c2v_parallelIn_304(c2v_in4[30]),
	.c2v_parallelIn_305(c2v_in5[30]),
	.c2v_parallelIn_310(c2v_in0[31]),
	.c2v_parallelIn_311(c2v_in1[31]),
	.c2v_parallelIn_312(c2v_in2[31]),
	.c2v_parallelIn_313(c2v_in3[31]),
	.c2v_parallelIn_314(c2v_in4[31]),
	.c2v_parallelIn_315(c2v_in5[31]),
	.c2v_parallelIn_320(c2v_in0[32]),
	.c2v_parallelIn_321(c2v_in1[32]),
	.c2v_parallelIn_322(c2v_in2[32]),
	.c2v_parallelIn_323(c2v_in3[32]),
	.c2v_parallelIn_324(c2v_in4[32]),
	.c2v_parallelIn_325(c2v_in5[32]),
	.c2v_parallelIn_330(c2v_in0[33]),
	.c2v_parallelIn_331(c2v_in1[33]),
	.c2v_parallelIn_332(c2v_in2[33]),
	.c2v_parallelIn_333(c2v_in3[33]),
	.c2v_parallelIn_334(c2v_in4[33]),
	.c2v_parallelIn_335(c2v_in5[33]),
	.c2v_parallelIn_340(c2v_in0[34]),
	.c2v_parallelIn_341(c2v_in1[34]),
	.c2v_parallelIn_342(c2v_in2[34]),
	.c2v_parallelIn_343(c2v_in3[34]),
	.c2v_parallelIn_344(c2v_in4[34]),
	.c2v_parallelIn_345(c2v_in5[34]),
	.c2v_parallelIn_350(c2v_in0[35]),
	.c2v_parallelIn_351(c2v_in1[35]),
	.c2v_parallelIn_352(c2v_in2[35]),
	.c2v_parallelIn_353(c2v_in3[35]),
	.c2v_parallelIn_354(c2v_in4[35]),
	.c2v_parallelIn_355(c2v_in5[35]),
	.c2v_parallelIn_360(c2v_in0[36]),
	.c2v_parallelIn_361(c2v_in1[36]),
	.c2v_parallelIn_362(c2v_in2[36]),
	.c2v_parallelIn_363(c2v_in3[36]),
	.c2v_parallelIn_364(c2v_in4[36]),
	.c2v_parallelIn_365(c2v_in5[36]),
	.c2v_parallelIn_370(c2v_in0[37]),
	.c2v_parallelIn_371(c2v_in1[37]),
	.c2v_parallelIn_372(c2v_in2[37]),
	.c2v_parallelIn_373(c2v_in3[37]),
	.c2v_parallelIn_374(c2v_in4[37]),
	.c2v_parallelIn_375(c2v_in5[37]),
	.c2v_parallelIn_380(c2v_in0[38]),
	.c2v_parallelIn_381(c2v_in1[38]),
	.c2v_parallelIn_382(c2v_in2[38]),
	.c2v_parallelIn_383(c2v_in3[38]),
	.c2v_parallelIn_384(c2v_in4[38]),
	.c2v_parallelIn_385(c2v_in5[38]),
	.c2v_parallelIn_390(c2v_in0[39]),
	.c2v_parallelIn_391(c2v_in1[39]),
	.c2v_parallelIn_392(c2v_in2[39]),
	.c2v_parallelIn_393(c2v_in3[39]),
	.c2v_parallelIn_394(c2v_in4[39]),
	.c2v_parallelIn_395(c2v_in5[39]),
	.c2v_parallelIn_400(c2v_in0[40]),
	.c2v_parallelIn_401(c2v_in1[40]),
	.c2v_parallelIn_402(c2v_in2[40]),
	.c2v_parallelIn_403(c2v_in3[40]),
	.c2v_parallelIn_404(c2v_in4[40]),
	.c2v_parallelIn_405(c2v_in5[40]),
	.c2v_parallelIn_410(c2v_in0[41]),
	.c2v_parallelIn_411(c2v_in1[41]),
	.c2v_parallelIn_412(c2v_in2[41]),
	.c2v_parallelIn_413(c2v_in3[41]),
	.c2v_parallelIn_414(c2v_in4[41]),
	.c2v_parallelIn_415(c2v_in5[41]),
	.c2v_parallelIn_420(c2v_in0[42]),
	.c2v_parallelIn_421(c2v_in1[42]),
	.c2v_parallelIn_422(c2v_in2[42]),
	.c2v_parallelIn_423(c2v_in3[42]),
	.c2v_parallelIn_424(c2v_in4[42]),
	.c2v_parallelIn_425(c2v_in5[42]),
	.c2v_parallelIn_430(c2v_in0[43]),
	.c2v_parallelIn_431(c2v_in1[43]),
	.c2v_parallelIn_432(c2v_in2[43]),
	.c2v_parallelIn_433(c2v_in3[43]),
	.c2v_parallelIn_434(c2v_in4[43]),
	.c2v_parallelIn_435(c2v_in5[43]),
	.c2v_parallelIn_440(c2v_in0[44]),
	.c2v_parallelIn_441(c2v_in1[44]),
	.c2v_parallelIn_442(c2v_in2[44]),
	.c2v_parallelIn_443(c2v_in3[44]),
	.c2v_parallelIn_444(c2v_in4[44]),
	.c2v_parallelIn_445(c2v_in5[44]),
	.c2v_parallelIn_450(c2v_in0[45]),
	.c2v_parallelIn_451(c2v_in1[45]),
	.c2v_parallelIn_452(c2v_in2[45]),
	.c2v_parallelIn_453(c2v_in3[45]),
	.c2v_parallelIn_454(c2v_in4[45]),
	.c2v_parallelIn_455(c2v_in5[45]),
	.c2v_parallelIn_460(c2v_in0[46]),
	.c2v_parallelIn_461(c2v_in1[46]),
	.c2v_parallelIn_462(c2v_in2[46]),
	.c2v_parallelIn_463(c2v_in3[46]),
	.c2v_parallelIn_464(c2v_in4[46]),
	.c2v_parallelIn_465(c2v_in5[46]),
	.c2v_parallelIn_470(c2v_in0[47]),
	.c2v_parallelIn_471(c2v_in1[47]),
	.c2v_parallelIn_472(c2v_in2[47]),
	.c2v_parallelIn_473(c2v_in3[47]),
	.c2v_parallelIn_474(c2v_in4[47]),
	.c2v_parallelIn_475(c2v_in5[47]),
	.c2v_parallelIn_480(c2v_in0[48]),
	.c2v_parallelIn_481(c2v_in1[48]),
	.c2v_parallelIn_482(c2v_in2[48]),
	.c2v_parallelIn_483(c2v_in3[48]),
	.c2v_parallelIn_484(c2v_in4[48]),
	.c2v_parallelIn_485(c2v_in5[48]),
	.c2v_parallelIn_490(c2v_in0[49]),
	.c2v_parallelIn_491(c2v_in1[49]),
	.c2v_parallelIn_492(c2v_in2[49]),
	.c2v_parallelIn_493(c2v_in3[49]),
	.c2v_parallelIn_494(c2v_in4[49]),
	.c2v_parallelIn_495(c2v_in5[49]),
	.c2v_parallelIn_500(c2v_in0[50]),
	.c2v_parallelIn_501(c2v_in1[50]),
	.c2v_parallelIn_502(c2v_in2[50]),
	.c2v_parallelIn_503(c2v_in3[50]),
	.c2v_parallelIn_504(c2v_in4[50]),
	.c2v_parallelIn_505(c2v_in5[50]),
	.c2v_parallelIn_510(c2v_in0[51]),
	.c2v_parallelIn_511(c2v_in1[51]),
	.c2v_parallelIn_512(c2v_in2[51]),
	.c2v_parallelIn_513(c2v_in3[51]),
	.c2v_parallelIn_514(c2v_in4[51]),
	.c2v_parallelIn_515(c2v_in5[51]),
	.c2v_parallelIn_520(c2v_in0[52]),
	.c2v_parallelIn_521(c2v_in1[52]),
	.c2v_parallelIn_522(c2v_in2[52]),
	.c2v_parallelIn_523(c2v_in3[52]),
	.c2v_parallelIn_524(c2v_in4[52]),
	.c2v_parallelIn_525(c2v_in5[52]),
	.c2v_parallelIn_530(c2v_in0[53]),
	.c2v_parallelIn_531(c2v_in1[53]),
	.c2v_parallelIn_532(c2v_in2[53]),
	.c2v_parallelIn_533(c2v_in3[53]),
	.c2v_parallelIn_534(c2v_in4[53]),
	.c2v_parallelIn_535(c2v_in5[53]),
	.c2v_parallelIn_540(c2v_in0[54]),
	.c2v_parallelIn_541(c2v_in1[54]),
	.c2v_parallelIn_542(c2v_in2[54]),
	.c2v_parallelIn_543(c2v_in3[54]),
	.c2v_parallelIn_544(c2v_in4[54]),
	.c2v_parallelIn_545(c2v_in5[54]),
	.c2v_parallelIn_550(c2v_in0[55]),
	.c2v_parallelIn_551(c2v_in1[55]),
	.c2v_parallelIn_552(c2v_in2[55]),
	.c2v_parallelIn_553(c2v_in3[55]),
	.c2v_parallelIn_554(c2v_in4[55]),
	.c2v_parallelIn_555(c2v_in5[55]),
	.c2v_parallelIn_560(c2v_in0[56]),
	.c2v_parallelIn_561(c2v_in1[56]),
	.c2v_parallelIn_562(c2v_in2[56]),
	.c2v_parallelIn_563(c2v_in3[56]),
	.c2v_parallelIn_564(c2v_in4[56]),
	.c2v_parallelIn_565(c2v_in5[56]),
	.c2v_parallelIn_570(c2v_in0[57]),
	.c2v_parallelIn_571(c2v_in1[57]),
	.c2v_parallelIn_572(c2v_in2[57]),
	.c2v_parallelIn_573(c2v_in3[57]),
	.c2v_parallelIn_574(c2v_in4[57]),
	.c2v_parallelIn_575(c2v_in5[57]),
	.c2v_parallelIn_580(c2v_in0[58]),
	.c2v_parallelIn_581(c2v_in1[58]),
	.c2v_parallelIn_582(c2v_in2[58]),
	.c2v_parallelIn_583(c2v_in3[58]),
	.c2v_parallelIn_584(c2v_in4[58]),
	.c2v_parallelIn_585(c2v_in5[58]),
	.c2v_parallelIn_590(c2v_in0[59]),
	.c2v_parallelIn_591(c2v_in1[59]),
	.c2v_parallelIn_592(c2v_in2[59]),
	.c2v_parallelIn_593(c2v_in3[59]),
	.c2v_parallelIn_594(c2v_in4[59]),
	.c2v_parallelIn_595(c2v_in5[59]),
	.c2v_parallelIn_600(c2v_in0[60]),
	.c2v_parallelIn_601(c2v_in1[60]),
	.c2v_parallelIn_602(c2v_in2[60]),
	.c2v_parallelIn_603(c2v_in3[60]),
	.c2v_parallelIn_604(c2v_in4[60]),
	.c2v_parallelIn_605(c2v_in5[60]),
	.c2v_parallelIn_610(c2v_in0[61]),
	.c2v_parallelIn_611(c2v_in1[61]),
	.c2v_parallelIn_612(c2v_in2[61]),
	.c2v_parallelIn_613(c2v_in3[61]),
	.c2v_parallelIn_614(c2v_in4[61]),
	.c2v_parallelIn_615(c2v_in5[61]),
	.c2v_parallelIn_620(c2v_in0[62]),
	.c2v_parallelIn_621(c2v_in1[62]),
	.c2v_parallelIn_622(c2v_in2[62]),
	.c2v_parallelIn_623(c2v_in3[62]),
	.c2v_parallelIn_624(c2v_in4[62]),
	.c2v_parallelIn_625(c2v_in5[62]),
	.c2v_parallelIn_630(c2v_in0[63]),
	.c2v_parallelIn_631(c2v_in1[63]),
	.c2v_parallelIn_632(c2v_in2[63]),
	.c2v_parallelIn_633(c2v_in3[63]),
	.c2v_parallelIn_634(c2v_in4[63]),
	.c2v_parallelIn_635(c2v_in5[63]),
	.c2v_parallelIn_640(c2v_in0[64]),
	.c2v_parallelIn_641(c2v_in1[64]),
	.c2v_parallelIn_642(c2v_in2[64]),
	.c2v_parallelIn_643(c2v_in3[64]),
	.c2v_parallelIn_644(c2v_in4[64]),
	.c2v_parallelIn_645(c2v_in5[64]),
	.c2v_parallelIn_650(c2v_in0[65]),
	.c2v_parallelIn_651(c2v_in1[65]),
	.c2v_parallelIn_652(c2v_in2[65]),
	.c2v_parallelIn_653(c2v_in3[65]),
	.c2v_parallelIn_654(c2v_in4[65]),
	.c2v_parallelIn_655(c2v_in5[65]),
	.c2v_parallelIn_660(c2v_in0[66]),
	.c2v_parallelIn_661(c2v_in1[66]),
	.c2v_parallelIn_662(c2v_in2[66]),
	.c2v_parallelIn_663(c2v_in3[66]),
	.c2v_parallelIn_664(c2v_in4[66]),
	.c2v_parallelIn_665(c2v_in5[66]),
	.c2v_parallelIn_670(c2v_in0[67]),
	.c2v_parallelIn_671(c2v_in1[67]),
	.c2v_parallelIn_672(c2v_in2[67]),
	.c2v_parallelIn_673(c2v_in3[67]),
	.c2v_parallelIn_674(c2v_in4[67]),
	.c2v_parallelIn_675(c2v_in5[67]),
	.c2v_parallelIn_680(c2v_in0[68]),
	.c2v_parallelIn_681(c2v_in1[68]),
	.c2v_parallelIn_682(c2v_in2[68]),
	.c2v_parallelIn_683(c2v_in3[68]),
	.c2v_parallelIn_684(c2v_in4[68]),
	.c2v_parallelIn_685(c2v_in5[68]),
	.c2v_parallelIn_690(c2v_in0[69]),
	.c2v_parallelIn_691(c2v_in1[69]),
	.c2v_parallelIn_692(c2v_in2[69]),
	.c2v_parallelIn_693(c2v_in3[69]),
	.c2v_parallelIn_694(c2v_in4[69]),
	.c2v_parallelIn_695(c2v_in5[69]),
	.c2v_parallelIn_700(c2v_in0[70]),
	.c2v_parallelIn_701(c2v_in1[70]),
	.c2v_parallelIn_702(c2v_in2[70]),
	.c2v_parallelIn_703(c2v_in3[70]),
	.c2v_parallelIn_704(c2v_in4[70]),
	.c2v_parallelIn_705(c2v_in5[70]),
	.c2v_parallelIn_710(c2v_in0[71]),
	.c2v_parallelIn_711(c2v_in1[71]),
	.c2v_parallelIn_712(c2v_in2[71]),
	.c2v_parallelIn_713(c2v_in3[71]),
	.c2v_parallelIn_714(c2v_in4[71]),
	.c2v_parallelIn_715(c2v_in5[71]),
	.c2v_parallelIn_720(c2v_in0[72]),
	.c2v_parallelIn_721(c2v_in1[72]),
	.c2v_parallelIn_722(c2v_in2[72]),
	.c2v_parallelIn_723(c2v_in3[72]),
	.c2v_parallelIn_724(c2v_in4[72]),
	.c2v_parallelIn_725(c2v_in5[72]),
	.c2v_parallelIn_730(c2v_in0[73]),
	.c2v_parallelIn_731(c2v_in1[73]),
	.c2v_parallelIn_732(c2v_in2[73]),
	.c2v_parallelIn_733(c2v_in3[73]),
	.c2v_parallelIn_734(c2v_in4[73]),
	.c2v_parallelIn_735(c2v_in5[73]),
	.c2v_parallelIn_740(c2v_in0[74]),
	.c2v_parallelIn_741(c2v_in1[74]),
	.c2v_parallelIn_742(c2v_in2[74]),
	.c2v_parallelIn_743(c2v_in3[74]),
	.c2v_parallelIn_744(c2v_in4[74]),
	.c2v_parallelIn_745(c2v_in5[74]),
	.c2v_parallelIn_750(c2v_in0[75]),
	.c2v_parallelIn_751(c2v_in1[75]),
	.c2v_parallelIn_752(c2v_in2[75]),
	.c2v_parallelIn_753(c2v_in3[75]),
	.c2v_parallelIn_754(c2v_in4[75]),
	.c2v_parallelIn_755(c2v_in5[75]),
	.c2v_parallelIn_760(c2v_in0[76]),
	.c2v_parallelIn_761(c2v_in1[76]),
	.c2v_parallelIn_762(c2v_in2[76]),
	.c2v_parallelIn_763(c2v_in3[76]),
	.c2v_parallelIn_764(c2v_in4[76]),
	.c2v_parallelIn_765(c2v_in5[76]),
	.c2v_parallelIn_770(c2v_in0[77]),
	.c2v_parallelIn_771(c2v_in1[77]),
	.c2v_parallelIn_772(c2v_in2[77]),
	.c2v_parallelIn_773(c2v_in3[77]),
	.c2v_parallelIn_774(c2v_in4[77]),
	.c2v_parallelIn_775(c2v_in5[77]),
	.c2v_parallelIn_780(c2v_in0[78]),
	.c2v_parallelIn_781(c2v_in1[78]),
	.c2v_parallelIn_782(c2v_in2[78]),
	.c2v_parallelIn_783(c2v_in3[78]),
	.c2v_parallelIn_784(c2v_in4[78]),
	.c2v_parallelIn_785(c2v_in5[78]),
	.c2v_parallelIn_790(c2v_in0[79]),
	.c2v_parallelIn_791(c2v_in1[79]),
	.c2v_parallelIn_792(c2v_in2[79]),
	.c2v_parallelIn_793(c2v_in3[79]),
	.c2v_parallelIn_794(c2v_in4[79]),
	.c2v_parallelIn_795(c2v_in5[79]),
	.c2v_parallelIn_800(c2v_in0[80]),
	.c2v_parallelIn_801(c2v_in1[80]),
	.c2v_parallelIn_802(c2v_in2[80]),
	.c2v_parallelIn_803(c2v_in3[80]),
	.c2v_parallelIn_804(c2v_in4[80]),
	.c2v_parallelIn_805(c2v_in5[80]),
	.c2v_parallelIn_810(c2v_in0[81]),
	.c2v_parallelIn_811(c2v_in1[81]),
	.c2v_parallelIn_812(c2v_in2[81]),
	.c2v_parallelIn_813(c2v_in3[81]),
	.c2v_parallelIn_814(c2v_in4[81]),
	.c2v_parallelIn_815(c2v_in5[81]),
	.c2v_parallelIn_820(c2v_in0[82]),
	.c2v_parallelIn_821(c2v_in1[82]),
	.c2v_parallelIn_822(c2v_in2[82]),
	.c2v_parallelIn_823(c2v_in3[82]),
	.c2v_parallelIn_824(c2v_in4[82]),
	.c2v_parallelIn_825(c2v_in5[82]),
	.c2v_parallelIn_830(c2v_in0[83]),
	.c2v_parallelIn_831(c2v_in1[83]),
	.c2v_parallelIn_832(c2v_in2[83]),
	.c2v_parallelIn_833(c2v_in3[83]),
	.c2v_parallelIn_834(c2v_in4[83]),
	.c2v_parallelIn_835(c2v_in5[83]),
	.c2v_parallelIn_840(c2v_in0[84]),
	.c2v_parallelIn_841(c2v_in1[84]),
	.c2v_parallelIn_842(c2v_in2[84]),
	.c2v_parallelIn_843(c2v_in3[84]),
	.c2v_parallelIn_844(c2v_in4[84]),
	.c2v_parallelIn_845(c2v_in5[84]),
	.c2v_parallelIn_850(c2v_in0[85]),
	.c2v_parallelIn_851(c2v_in1[85]),
	.c2v_parallelIn_852(c2v_in2[85]),
	.c2v_parallelIn_853(c2v_in3[85]),
	.c2v_parallelIn_854(c2v_in4[85]),
	.c2v_parallelIn_855(c2v_in5[85]),
	.c2v_parallelIn_860(c2v_in0[86]),
	.c2v_parallelIn_861(c2v_in1[86]),
	.c2v_parallelIn_862(c2v_in2[86]),
	.c2v_parallelIn_863(c2v_in3[86]),
	.c2v_parallelIn_864(c2v_in4[86]),
	.c2v_parallelIn_865(c2v_in5[86]),
	.c2v_parallelIn_870(c2v_in0[87]),
	.c2v_parallelIn_871(c2v_in1[87]),
	.c2v_parallelIn_872(c2v_in2[87]),
	.c2v_parallelIn_873(c2v_in3[87]),
	.c2v_parallelIn_874(c2v_in4[87]),
	.c2v_parallelIn_875(c2v_in5[87]),
	.c2v_parallelIn_880(c2v_in0[88]),
	.c2v_parallelIn_881(c2v_in1[88]),
	.c2v_parallelIn_882(c2v_in2[88]),
	.c2v_parallelIn_883(c2v_in3[88]),
	.c2v_parallelIn_884(c2v_in4[88]),
	.c2v_parallelIn_885(c2v_in5[88]),
	.c2v_parallelIn_890(c2v_in0[89]),
	.c2v_parallelIn_891(c2v_in1[89]),
	.c2v_parallelIn_892(c2v_in2[89]),
	.c2v_parallelIn_893(c2v_in3[89]),
	.c2v_parallelIn_894(c2v_in4[89]),
	.c2v_parallelIn_895(c2v_in5[89]),
	.c2v_parallelIn_900(c2v_in0[90]),
	.c2v_parallelIn_901(c2v_in1[90]),
	.c2v_parallelIn_902(c2v_in2[90]),
	.c2v_parallelIn_903(c2v_in3[90]),
	.c2v_parallelIn_904(c2v_in4[90]),
	.c2v_parallelIn_905(c2v_in5[90]),
	.c2v_parallelIn_910(c2v_in0[91]),
	.c2v_parallelIn_911(c2v_in1[91]),
	.c2v_parallelIn_912(c2v_in2[91]),
	.c2v_parallelIn_913(c2v_in3[91]),
	.c2v_parallelIn_914(c2v_in4[91]),
	.c2v_parallelIn_915(c2v_in5[91]),
	.c2v_parallelIn_920(c2v_in0[92]),
	.c2v_parallelIn_921(c2v_in1[92]),
	.c2v_parallelIn_922(c2v_in2[92]),
	.c2v_parallelIn_923(c2v_in3[92]),
	.c2v_parallelIn_924(c2v_in4[92]),
	.c2v_parallelIn_925(c2v_in5[92]),
	.c2v_parallelIn_930(c2v_in0[93]),
	.c2v_parallelIn_931(c2v_in1[93]),
	.c2v_parallelIn_932(c2v_in2[93]),
	.c2v_parallelIn_933(c2v_in3[93]),
	.c2v_parallelIn_934(c2v_in4[93]),
	.c2v_parallelIn_935(c2v_in5[93]),
	.c2v_parallelIn_940(c2v_in0[94]),
	.c2v_parallelIn_941(c2v_in1[94]),
	.c2v_parallelIn_942(c2v_in2[94]),
	.c2v_parallelIn_943(c2v_in3[94]),
	.c2v_parallelIn_944(c2v_in4[94]),
	.c2v_parallelIn_945(c2v_in5[94]),
	.c2v_parallelIn_950(c2v_in0[95]),
	.c2v_parallelIn_951(c2v_in1[95]),
	.c2v_parallelIn_952(c2v_in2[95]),
	.c2v_parallelIn_953(c2v_in3[95]),
	.c2v_parallelIn_954(c2v_in4[95]),
	.c2v_parallelIn_955(c2v_in5[95]),
	.c2v_parallelIn_960(c2v_in0[96]),
	.c2v_parallelIn_961(c2v_in1[96]),
	.c2v_parallelIn_962(c2v_in2[96]),
	.c2v_parallelIn_963(c2v_in3[96]),
	.c2v_parallelIn_964(c2v_in4[96]),
	.c2v_parallelIn_965(c2v_in5[96]),
	.c2v_parallelIn_970(c2v_in0[97]),
	.c2v_parallelIn_971(c2v_in1[97]),
	.c2v_parallelIn_972(c2v_in2[97]),
	.c2v_parallelIn_973(c2v_in3[97]),
	.c2v_parallelIn_974(c2v_in4[97]),
	.c2v_parallelIn_975(c2v_in5[97]),
	.c2v_parallelIn_980(c2v_in0[98]),
	.c2v_parallelIn_981(c2v_in1[98]),
	.c2v_parallelIn_982(c2v_in2[98]),
	.c2v_parallelIn_983(c2v_in3[98]),
	.c2v_parallelIn_984(c2v_in4[98]),
	.c2v_parallelIn_985(c2v_in5[98]),
	.c2v_parallelIn_990(c2v_in0[99]),
	.c2v_parallelIn_991(c2v_in1[99]),
	.c2v_parallelIn_992(c2v_in2[99]),
	.c2v_parallelIn_993(c2v_in3[99]),
	.c2v_parallelIn_994(c2v_in4[99]),
	.c2v_parallelIn_995(c2v_in5[99]),
	.c2v_parallelIn_1000(c2v_in0[100]),
	.c2v_parallelIn_1001(c2v_in1[100]),
	.c2v_parallelIn_1002(c2v_in2[100]),
	.c2v_parallelIn_1003(c2v_in3[100]),
	.c2v_parallelIn_1004(c2v_in4[100]),
	.c2v_parallelIn_1005(c2v_in5[100]),
	.c2v_parallelIn_1010(c2v_in0[101]),
	.c2v_parallelIn_1011(c2v_in1[101]),
	.c2v_parallelIn_1012(c2v_in2[101]),
	.c2v_parallelIn_1013(c2v_in3[101]),
	.c2v_parallelIn_1014(c2v_in4[101]),
	.c2v_parallelIn_1015(c2v_in5[101]),
	
	.v2c_parallelIn_00(v2c_in0[0]),
	.v2c_parallelIn_01(v2c_in1[0]),
	.v2c_parallelIn_02(v2c_in2[0]),
	.v2c_parallelIn_10(v2c_in0[1]),
	.v2c_parallelIn_11(v2c_in1[1]),
	.v2c_parallelIn_12(v2c_in2[1]),
	.v2c_parallelIn_20(v2c_in0[2]),
	.v2c_parallelIn_21(v2c_in1[2]),
	.v2c_parallelIn_22(v2c_in2[2]),
	.v2c_parallelIn_30(v2c_in0[3]),
	.v2c_parallelIn_31(v2c_in1[3]),
	.v2c_parallelIn_32(v2c_in2[3]),
	.v2c_parallelIn_40(v2c_in0[4]),
	.v2c_parallelIn_41(v2c_in1[4]),
	.v2c_parallelIn_42(v2c_in2[4]),
	.v2c_parallelIn_50(v2c_in0[5]),
	.v2c_parallelIn_51(v2c_in1[5]),
	.v2c_parallelIn_52(v2c_in2[5]),
	.v2c_parallelIn_60(v2c_in0[6]),
	.v2c_parallelIn_61(v2c_in1[6]),
	.v2c_parallelIn_62(v2c_in2[6]),
	.v2c_parallelIn_70(v2c_in0[7]),
	.v2c_parallelIn_71(v2c_in1[7]),
	.v2c_parallelIn_72(v2c_in2[7]),
	.v2c_parallelIn_80(v2c_in0[8]),
	.v2c_parallelIn_81(v2c_in1[8]),
	.v2c_parallelIn_82(v2c_in2[8]),
	.v2c_parallelIn_90(v2c_in0[9]),
	.v2c_parallelIn_91(v2c_in1[9]),
	.v2c_parallelIn_92(v2c_in2[9]),
	.v2c_parallelIn_100(v2c_in0[10]),
	.v2c_parallelIn_101(v2c_in1[10]),
	.v2c_parallelIn_102(v2c_in2[10]),
	.v2c_parallelIn_110(v2c_in0[11]),
	.v2c_parallelIn_111(v2c_in1[11]),
	.v2c_parallelIn_112(v2c_in2[11]),
	.v2c_parallelIn_120(v2c_in0[12]),
	.v2c_parallelIn_121(v2c_in1[12]),
	.v2c_parallelIn_122(v2c_in2[12]),
	.v2c_parallelIn_130(v2c_in0[13]),
	.v2c_parallelIn_131(v2c_in1[13]),
	.v2c_parallelIn_132(v2c_in2[13]),
	.v2c_parallelIn_140(v2c_in0[14]),
	.v2c_parallelIn_141(v2c_in1[14]),
	.v2c_parallelIn_142(v2c_in2[14]),
	.v2c_parallelIn_150(v2c_in0[15]),
	.v2c_parallelIn_151(v2c_in1[15]),
	.v2c_parallelIn_152(v2c_in2[15]),
	.v2c_parallelIn_160(v2c_in0[16]),
	.v2c_parallelIn_161(v2c_in1[16]),
	.v2c_parallelIn_162(v2c_in2[16]),
	.v2c_parallelIn_170(v2c_in0[17]),
	.v2c_parallelIn_171(v2c_in1[17]),
	.v2c_parallelIn_172(v2c_in2[17]),
	.v2c_parallelIn_180(v2c_in0[18]),
	.v2c_parallelIn_181(v2c_in1[18]),
	.v2c_parallelIn_182(v2c_in2[18]),
	.v2c_parallelIn_190(v2c_in0[19]),
	.v2c_parallelIn_191(v2c_in1[19]),
	.v2c_parallelIn_192(v2c_in2[19]),
	.v2c_parallelIn_200(v2c_in0[20]),
	.v2c_parallelIn_201(v2c_in1[20]),
	.v2c_parallelIn_202(v2c_in2[20]),
	.v2c_parallelIn_210(v2c_in0[21]),
	.v2c_parallelIn_211(v2c_in1[21]),
	.v2c_parallelIn_212(v2c_in2[21]),
	.v2c_parallelIn_220(v2c_in0[22]),
	.v2c_parallelIn_221(v2c_in1[22]),
	.v2c_parallelIn_222(v2c_in2[22]),
	.v2c_parallelIn_230(v2c_in0[23]),
	.v2c_parallelIn_231(v2c_in1[23]),
	.v2c_parallelIn_232(v2c_in2[23]),
	.v2c_parallelIn_240(v2c_in0[24]),
	.v2c_parallelIn_241(v2c_in1[24]),
	.v2c_parallelIn_242(v2c_in2[24]),
	.v2c_parallelIn_250(v2c_in0[25]),
	.v2c_parallelIn_251(v2c_in1[25]),
	.v2c_parallelIn_252(v2c_in2[25]),
	.v2c_parallelIn_260(v2c_in0[26]),
	.v2c_parallelIn_261(v2c_in1[26]),
	.v2c_parallelIn_262(v2c_in2[26]),
	.v2c_parallelIn_270(v2c_in0[27]),
	.v2c_parallelIn_271(v2c_in1[27]),
	.v2c_parallelIn_272(v2c_in2[27]),
	.v2c_parallelIn_280(v2c_in0[28]),
	.v2c_parallelIn_281(v2c_in1[28]),
	.v2c_parallelIn_282(v2c_in2[28]),
	.v2c_parallelIn_290(v2c_in0[29]),
	.v2c_parallelIn_291(v2c_in1[29]),
	.v2c_parallelIn_292(v2c_in2[29]),
	.v2c_parallelIn_300(v2c_in0[30]),
	.v2c_parallelIn_301(v2c_in1[30]),
	.v2c_parallelIn_302(v2c_in2[30]),
	.v2c_parallelIn_310(v2c_in0[31]),
	.v2c_parallelIn_311(v2c_in1[31]),
	.v2c_parallelIn_312(v2c_in2[31]),
	.v2c_parallelIn_320(v2c_in0[32]),
	.v2c_parallelIn_321(v2c_in1[32]),
	.v2c_parallelIn_322(v2c_in2[32]),
	.v2c_parallelIn_330(v2c_in0[33]),
	.v2c_parallelIn_331(v2c_in1[33]),
	.v2c_parallelIn_332(v2c_in2[33]),
	.v2c_parallelIn_340(v2c_in0[34]),
	.v2c_parallelIn_341(v2c_in1[34]),
	.v2c_parallelIn_342(v2c_in2[34]),
	.v2c_parallelIn_350(v2c_in0[35]),
	.v2c_parallelIn_351(v2c_in1[35]),
	.v2c_parallelIn_352(v2c_in2[35]),
	.v2c_parallelIn_360(v2c_in0[36]),
	.v2c_parallelIn_361(v2c_in1[36]),
	.v2c_parallelIn_362(v2c_in2[36]),
	.v2c_parallelIn_370(v2c_in0[37]),
	.v2c_parallelIn_371(v2c_in1[37]),
	.v2c_parallelIn_372(v2c_in2[37]),
	.v2c_parallelIn_380(v2c_in0[38]),
	.v2c_parallelIn_381(v2c_in1[38]),
	.v2c_parallelIn_382(v2c_in2[38]),
	.v2c_parallelIn_390(v2c_in0[39]),
	.v2c_parallelIn_391(v2c_in1[39]),
	.v2c_parallelIn_392(v2c_in2[39]),
	.v2c_parallelIn_400(v2c_in0[40]),
	.v2c_parallelIn_401(v2c_in1[40]),
	.v2c_parallelIn_402(v2c_in2[40]),
	.v2c_parallelIn_410(v2c_in0[41]),
	.v2c_parallelIn_411(v2c_in1[41]),
	.v2c_parallelIn_412(v2c_in2[41]),
	.v2c_parallelIn_420(v2c_in0[42]),
	.v2c_parallelIn_421(v2c_in1[42]),
	.v2c_parallelIn_422(v2c_in2[42]),
	.v2c_parallelIn_430(v2c_in0[43]),
	.v2c_parallelIn_431(v2c_in1[43]),
	.v2c_parallelIn_432(v2c_in2[43]),
	.v2c_parallelIn_440(v2c_in0[44]),
	.v2c_parallelIn_441(v2c_in1[44]),
	.v2c_parallelIn_442(v2c_in2[44]),
	.v2c_parallelIn_450(v2c_in0[45]),
	.v2c_parallelIn_451(v2c_in1[45]),
	.v2c_parallelIn_452(v2c_in2[45]),
	.v2c_parallelIn_460(v2c_in0[46]),
	.v2c_parallelIn_461(v2c_in1[46]),
	.v2c_parallelIn_462(v2c_in2[46]),
	.v2c_parallelIn_470(v2c_in0[47]),
	.v2c_parallelIn_471(v2c_in1[47]),
	.v2c_parallelIn_472(v2c_in2[47]),
	.v2c_parallelIn_480(v2c_in0[48]),
	.v2c_parallelIn_481(v2c_in1[48]),
	.v2c_parallelIn_482(v2c_in2[48]),
	.v2c_parallelIn_490(v2c_in0[49]),
	.v2c_parallelIn_491(v2c_in1[49]),
	.v2c_parallelIn_492(v2c_in2[49]),
	.v2c_parallelIn_500(v2c_in0[50]),
	.v2c_parallelIn_501(v2c_in1[50]),
	.v2c_parallelIn_502(v2c_in2[50]),
	.v2c_parallelIn_510(v2c_in0[51]),
	.v2c_parallelIn_511(v2c_in1[51]),
	.v2c_parallelIn_512(v2c_in2[51]),
	.v2c_parallelIn_520(v2c_in0[52]),
	.v2c_parallelIn_521(v2c_in1[52]),
	.v2c_parallelIn_522(v2c_in2[52]),
	.v2c_parallelIn_530(v2c_in0[53]),
	.v2c_parallelIn_531(v2c_in1[53]),
	.v2c_parallelIn_532(v2c_in2[53]),
	.v2c_parallelIn_540(v2c_in0[54]),
	.v2c_parallelIn_541(v2c_in1[54]),
	.v2c_parallelIn_542(v2c_in2[54]),
	.v2c_parallelIn_550(v2c_in0[55]),
	.v2c_parallelIn_551(v2c_in1[55]),
	.v2c_parallelIn_552(v2c_in2[55]),
	.v2c_parallelIn_560(v2c_in0[56]),
	.v2c_parallelIn_561(v2c_in1[56]),
	.v2c_parallelIn_562(v2c_in2[56]),
	.v2c_parallelIn_570(v2c_in0[57]),
	.v2c_parallelIn_571(v2c_in1[57]),
	.v2c_parallelIn_572(v2c_in2[57]),
	.v2c_parallelIn_580(v2c_in0[58]),
	.v2c_parallelIn_581(v2c_in1[58]),
	.v2c_parallelIn_582(v2c_in2[58]),
	.v2c_parallelIn_590(v2c_in0[59]),
	.v2c_parallelIn_591(v2c_in1[59]),
	.v2c_parallelIn_592(v2c_in2[59]),
	.v2c_parallelIn_600(v2c_in0[60]),
	.v2c_parallelIn_601(v2c_in1[60]),
	.v2c_parallelIn_602(v2c_in2[60]),
	.v2c_parallelIn_610(v2c_in0[61]),
	.v2c_parallelIn_611(v2c_in1[61]),
	.v2c_parallelIn_612(v2c_in2[61]),
	.v2c_parallelIn_620(v2c_in0[62]),
	.v2c_parallelIn_621(v2c_in1[62]),
	.v2c_parallelIn_622(v2c_in2[62]),
	.v2c_parallelIn_630(v2c_in0[63]),
	.v2c_parallelIn_631(v2c_in1[63]),
	.v2c_parallelIn_632(v2c_in2[63]),
	.v2c_parallelIn_640(v2c_in0[64]),
	.v2c_parallelIn_641(v2c_in1[64]),
	.v2c_parallelIn_642(v2c_in2[64]),
	.v2c_parallelIn_650(v2c_in0[65]),
	.v2c_parallelIn_651(v2c_in1[65]),
	.v2c_parallelIn_652(v2c_in2[65]),
	.v2c_parallelIn_660(v2c_in0[66]),
	.v2c_parallelIn_661(v2c_in1[66]),
	.v2c_parallelIn_662(v2c_in2[66]),
	.v2c_parallelIn_670(v2c_in0[67]),
	.v2c_parallelIn_671(v2c_in1[67]),
	.v2c_parallelIn_672(v2c_in2[67]),
	.v2c_parallelIn_680(v2c_in0[68]),
	.v2c_parallelIn_681(v2c_in1[68]),
	.v2c_parallelIn_682(v2c_in2[68]),
	.v2c_parallelIn_690(v2c_in0[69]),
	.v2c_parallelIn_691(v2c_in1[69]),
	.v2c_parallelIn_692(v2c_in2[69]),
	.v2c_parallelIn_700(v2c_in0[70]),
	.v2c_parallelIn_701(v2c_in1[70]),
	.v2c_parallelIn_702(v2c_in2[70]),
	.v2c_parallelIn_710(v2c_in0[71]),
	.v2c_parallelIn_711(v2c_in1[71]),
	.v2c_parallelIn_712(v2c_in2[71]),
	.v2c_parallelIn_720(v2c_in0[72]),
	.v2c_parallelIn_721(v2c_in1[72]),
	.v2c_parallelIn_722(v2c_in2[72]),
	.v2c_parallelIn_730(v2c_in0[73]),
	.v2c_parallelIn_731(v2c_in1[73]),
	.v2c_parallelIn_732(v2c_in2[73]),
	.v2c_parallelIn_740(v2c_in0[74]),
	.v2c_parallelIn_741(v2c_in1[74]),
	.v2c_parallelIn_742(v2c_in2[74]),
	.v2c_parallelIn_750(v2c_in0[75]),
	.v2c_parallelIn_751(v2c_in1[75]),
	.v2c_parallelIn_752(v2c_in2[75]),
	.v2c_parallelIn_760(v2c_in0[76]),
	.v2c_parallelIn_761(v2c_in1[76]),
	.v2c_parallelIn_762(v2c_in2[76]),
	.v2c_parallelIn_770(v2c_in0[77]),
	.v2c_parallelIn_771(v2c_in1[77]),
	.v2c_parallelIn_772(v2c_in2[77]),
	.v2c_parallelIn_780(v2c_in0[78]),
	.v2c_parallelIn_781(v2c_in1[78]),
	.v2c_parallelIn_782(v2c_in2[78]),
	.v2c_parallelIn_790(v2c_in0[79]),
	.v2c_parallelIn_791(v2c_in1[79]),
	.v2c_parallelIn_792(v2c_in2[79]),
	.v2c_parallelIn_800(v2c_in0[80]),
	.v2c_parallelIn_801(v2c_in1[80]),
	.v2c_parallelIn_802(v2c_in2[80]),
	.v2c_parallelIn_810(v2c_in0[81]),
	.v2c_parallelIn_811(v2c_in1[81]),
	.v2c_parallelIn_812(v2c_in2[81]),
	.v2c_parallelIn_820(v2c_in0[82]),
	.v2c_parallelIn_821(v2c_in1[82]),
	.v2c_parallelIn_822(v2c_in2[82]),
	.v2c_parallelIn_830(v2c_in0[83]),
	.v2c_parallelIn_831(v2c_in1[83]),
	.v2c_parallelIn_832(v2c_in2[83]),
	.v2c_parallelIn_840(v2c_in0[84]),
	.v2c_parallelIn_841(v2c_in1[84]),
	.v2c_parallelIn_842(v2c_in2[84]),
	.v2c_parallelIn_850(v2c_in0[85]),
	.v2c_parallelIn_851(v2c_in1[85]),
	.v2c_parallelIn_852(v2c_in2[85]),
	.v2c_parallelIn_860(v2c_in0[86]),
	.v2c_parallelIn_861(v2c_in1[86]),
	.v2c_parallelIn_862(v2c_in2[86]),
	.v2c_parallelIn_870(v2c_in0[87]),
	.v2c_parallelIn_871(v2c_in1[87]),
	.v2c_parallelIn_872(v2c_in2[87]),
	.v2c_parallelIn_880(v2c_in0[88]),
	.v2c_parallelIn_881(v2c_in1[88]),
	.v2c_parallelIn_882(v2c_in2[88]),
	.v2c_parallelIn_890(v2c_in0[89]),
	.v2c_parallelIn_891(v2c_in1[89]),
	.v2c_parallelIn_892(v2c_in2[89]),
	.v2c_parallelIn_900(v2c_in0[90]),
	.v2c_parallelIn_901(v2c_in1[90]),
	.v2c_parallelIn_902(v2c_in2[90]),
	.v2c_parallelIn_910(v2c_in0[91]),
	.v2c_parallelIn_911(v2c_in1[91]),
	.v2c_parallelIn_912(v2c_in2[91]),
	.v2c_parallelIn_920(v2c_in0[92]),
	.v2c_parallelIn_921(v2c_in1[92]),
	.v2c_parallelIn_922(v2c_in2[92]),
	.v2c_parallelIn_930(v2c_in0[93]),
	.v2c_parallelIn_931(v2c_in1[93]),
	.v2c_parallelIn_932(v2c_in2[93]),
	.v2c_parallelIn_940(v2c_in0[94]),
	.v2c_parallelIn_941(v2c_in1[94]),
	.v2c_parallelIn_942(v2c_in2[94]),
	.v2c_parallelIn_950(v2c_in0[95]),
	.v2c_parallelIn_951(v2c_in1[95]),
	.v2c_parallelIn_952(v2c_in2[95]),
	.v2c_parallelIn_960(v2c_in0[96]),
	.v2c_parallelIn_961(v2c_in1[96]),
	.v2c_parallelIn_962(v2c_in2[96]),
	.v2c_parallelIn_970(v2c_in0[97]),
	.v2c_parallelIn_971(v2c_in1[97]),
	.v2c_parallelIn_972(v2c_in2[97]),
	.v2c_parallelIn_980(v2c_in0[98]),
	.v2c_parallelIn_981(v2c_in1[98]),
	.v2c_parallelIn_982(v2c_in2[98]),
	.v2c_parallelIn_990(v2c_in0[99]),
	.v2c_parallelIn_991(v2c_in1[99]),
	.v2c_parallelIn_992(v2c_in2[99]),
	.v2c_parallelIn_1000(v2c_in0[100]),
	.v2c_parallelIn_1001(v2c_in1[100]),
	.v2c_parallelIn_1002(v2c_in2[100]),
	.v2c_parallelIn_1010(v2c_in0[101]),
	.v2c_parallelIn_1011(v2c_in1[101]),
	.v2c_parallelIn_1012(v2c_in2[101]),
	.v2c_parallelIn_1020(v2c_in0[102]),
	.v2c_parallelIn_1021(v2c_in1[102]),
	.v2c_parallelIn_1022(v2c_in2[102]),
	.v2c_parallelIn_1030(v2c_in0[103]),
	.v2c_parallelIn_1031(v2c_in1[103]),
	.v2c_parallelIn_1032(v2c_in2[103]),
	.v2c_parallelIn_1040(v2c_in0[104]),
	.v2c_parallelIn_1041(v2c_in1[104]),
	.v2c_parallelIn_1042(v2c_in2[104]),
	.v2c_parallelIn_1050(v2c_in0[105]),
	.v2c_parallelIn_1051(v2c_in1[105]),
	.v2c_parallelIn_1052(v2c_in2[105]),
	.v2c_parallelIn_1060(v2c_in0[106]),
	.v2c_parallelIn_1061(v2c_in1[106]),
	.v2c_parallelIn_1062(v2c_in2[106]),
	.v2c_parallelIn_1070(v2c_in0[107]),
	.v2c_parallelIn_1071(v2c_in1[107]),
	.v2c_parallelIn_1072(v2c_in2[107]),
	.v2c_parallelIn_1080(v2c_in0[108]),
	.v2c_parallelIn_1081(v2c_in1[108]),
	.v2c_parallelIn_1082(v2c_in2[108]),
	.v2c_parallelIn_1090(v2c_in0[109]),
	.v2c_parallelIn_1091(v2c_in1[109]),
	.v2c_parallelIn_1092(v2c_in2[109]),
	.v2c_parallelIn_1100(v2c_in0[110]),
	.v2c_parallelIn_1101(v2c_in1[110]),
	.v2c_parallelIn_1102(v2c_in2[110]),
	.v2c_parallelIn_1110(v2c_in0[111]),
	.v2c_parallelIn_1111(v2c_in1[111]),
	.v2c_parallelIn_1112(v2c_in2[111]),
	.v2c_parallelIn_1120(v2c_in0[112]),
	.v2c_parallelIn_1121(v2c_in1[112]),
	.v2c_parallelIn_1122(v2c_in2[112]),
	.v2c_parallelIn_1130(v2c_in0[113]),
	.v2c_parallelIn_1131(v2c_in1[113]),
	.v2c_parallelIn_1132(v2c_in2[113]),
	.v2c_parallelIn_1140(v2c_in0[114]),
	.v2c_parallelIn_1141(v2c_in1[114]),
	.v2c_parallelIn_1142(v2c_in2[114]),
	.v2c_parallelIn_1150(v2c_in0[115]),
	.v2c_parallelIn_1151(v2c_in1[115]),
	.v2c_parallelIn_1152(v2c_in2[115]),
	.v2c_parallelIn_1160(v2c_in0[116]),
	.v2c_parallelIn_1161(v2c_in1[116]),
	.v2c_parallelIn_1162(v2c_in2[116]),
	.v2c_parallelIn_1170(v2c_in0[117]),
	.v2c_parallelIn_1171(v2c_in1[117]),
	.v2c_parallelIn_1172(v2c_in2[117]),
	.v2c_parallelIn_1180(v2c_in0[118]),
	.v2c_parallelIn_1181(v2c_in1[118]),
	.v2c_parallelIn_1182(v2c_in2[118]),
	.v2c_parallelIn_1190(v2c_in0[119]),
	.v2c_parallelIn_1191(v2c_in1[119]),
	.v2c_parallelIn_1192(v2c_in2[119]),
	.v2c_parallelIn_1200(v2c_in0[120]),
	.v2c_parallelIn_1201(v2c_in1[120]),
	.v2c_parallelIn_1202(v2c_in2[120]),
	.v2c_parallelIn_1210(v2c_in0[121]),
	.v2c_parallelIn_1211(v2c_in1[121]),
	.v2c_parallelIn_1212(v2c_in2[121]),
	.v2c_parallelIn_1220(v2c_in0[122]),
	.v2c_parallelIn_1221(v2c_in1[122]),
	.v2c_parallelIn_1222(v2c_in2[122]),
	.v2c_parallelIn_1230(v2c_in0[123]),
	.v2c_parallelIn_1231(v2c_in1[123]),
	.v2c_parallelIn_1232(v2c_in2[123]),
	.v2c_parallelIn_1240(v2c_in0[124]),
	.v2c_parallelIn_1241(v2c_in1[124]),
	.v2c_parallelIn_1242(v2c_in2[124]),
	.v2c_parallelIn_1250(v2c_in0[125]),
	.v2c_parallelIn_1251(v2c_in1[125]),
	.v2c_parallelIn_1252(v2c_in2[125]),
	.v2c_parallelIn_1260(v2c_in0[126]),
	.v2c_parallelIn_1261(v2c_in1[126]),
	.v2c_parallelIn_1262(v2c_in2[126]),
	.v2c_parallelIn_1270(v2c_in0[127]),
	.v2c_parallelIn_1271(v2c_in1[127]),
	.v2c_parallelIn_1272(v2c_in2[127]),
	.v2c_parallelIn_1280(v2c_in0[128]),
	.v2c_parallelIn_1281(v2c_in1[128]),
	.v2c_parallelIn_1282(v2c_in2[128]),
	.v2c_parallelIn_1290(v2c_in0[129]),
	.v2c_parallelIn_1291(v2c_in1[129]),
	.v2c_parallelIn_1292(v2c_in2[129]),
	.v2c_parallelIn_1300(v2c_in0[130]),
	.v2c_parallelIn_1301(v2c_in1[130]),
	.v2c_parallelIn_1302(v2c_in2[130]),
	.v2c_parallelIn_1310(v2c_in0[131]),
	.v2c_parallelIn_1311(v2c_in1[131]),
	.v2c_parallelIn_1312(v2c_in2[131]),
	.v2c_parallelIn_1320(v2c_in0[132]),
	.v2c_parallelIn_1321(v2c_in1[132]),
	.v2c_parallelIn_1322(v2c_in2[132]),
	.v2c_parallelIn_1330(v2c_in0[133]),
	.v2c_parallelIn_1331(v2c_in1[133]),
	.v2c_parallelIn_1332(v2c_in2[133]),
	.v2c_parallelIn_1340(v2c_in0[134]),
	.v2c_parallelIn_1341(v2c_in1[134]),
	.v2c_parallelIn_1342(v2c_in2[134]),
	.v2c_parallelIn_1350(v2c_in0[135]),
	.v2c_parallelIn_1351(v2c_in1[135]),
	.v2c_parallelIn_1352(v2c_in2[135]),
	.v2c_parallelIn_1360(v2c_in0[136]),
	.v2c_parallelIn_1361(v2c_in1[136]),
	.v2c_parallelIn_1362(v2c_in2[136]),
	.v2c_parallelIn_1370(v2c_in0[137]),
	.v2c_parallelIn_1371(v2c_in1[137]),
	.v2c_parallelIn_1372(v2c_in2[137]),
	.v2c_parallelIn_1380(v2c_in0[138]),
	.v2c_parallelIn_1381(v2c_in1[138]),
	.v2c_parallelIn_1382(v2c_in2[138]),
	.v2c_parallelIn_1390(v2c_in0[139]),
	.v2c_parallelIn_1391(v2c_in1[139]),
	.v2c_parallelIn_1392(v2c_in2[139]),
	.v2c_parallelIn_1400(v2c_in0[140]),
	.v2c_parallelIn_1401(v2c_in1[140]),
	.v2c_parallelIn_1402(v2c_in2[140]),
	.v2c_parallelIn_1410(v2c_in0[141]),
	.v2c_parallelIn_1411(v2c_in1[141]),
	.v2c_parallelIn_1412(v2c_in2[141]),
	.v2c_parallelIn_1420(v2c_in0[142]),
	.v2c_parallelIn_1421(v2c_in1[142]),
	.v2c_parallelIn_1422(v2c_in2[142]),
	.v2c_parallelIn_1430(v2c_in0[143]),
	.v2c_parallelIn_1431(v2c_in1[143]),
	.v2c_parallelIn_1432(v2c_in2[143]),
	.v2c_parallelIn_1440(v2c_in0[144]),
	.v2c_parallelIn_1441(v2c_in1[144]),
	.v2c_parallelIn_1442(v2c_in2[144]),
	.v2c_parallelIn_1450(v2c_in0[145]),
	.v2c_parallelIn_1451(v2c_in1[145]),
	.v2c_parallelIn_1452(v2c_in2[145]),
	.v2c_parallelIn_1460(v2c_in0[146]),
	.v2c_parallelIn_1461(v2c_in1[146]),
	.v2c_parallelIn_1462(v2c_in2[146]),
	.v2c_parallelIn_1470(v2c_in0[147]),
	.v2c_parallelIn_1471(v2c_in1[147]),
	.v2c_parallelIn_1472(v2c_in2[147]),
	.v2c_parallelIn_1480(v2c_in0[148]),
	.v2c_parallelIn_1481(v2c_in1[148]),
	.v2c_parallelIn_1482(v2c_in2[148]),
	.v2c_parallelIn_1490(v2c_in0[149]),
	.v2c_parallelIn_1491(v2c_in1[149]),
	.v2c_parallelIn_1492(v2c_in2[149]),
	.v2c_parallelIn_1500(v2c_in0[150]),
	.v2c_parallelIn_1501(v2c_in1[150]),
	.v2c_parallelIn_1502(v2c_in2[150]),
	.v2c_parallelIn_1510(v2c_in0[151]),
	.v2c_parallelIn_1511(v2c_in1[151]),
	.v2c_parallelIn_1512(v2c_in2[151]),
	.v2c_parallelIn_1520(v2c_in0[152]),
	.v2c_parallelIn_1521(v2c_in1[152]),
	.v2c_parallelIn_1522(v2c_in2[152]),
	.v2c_parallelIn_1530(v2c_in0[153]),
	.v2c_parallelIn_1531(v2c_in1[153]),
	.v2c_parallelIn_1532(v2c_in2[153]),
	.v2c_parallelIn_1540(v2c_in0[154]),
	.v2c_parallelIn_1541(v2c_in1[154]),
	.v2c_parallelIn_1542(v2c_in2[154]),
	.v2c_parallelIn_1550(v2c_in0[155]),
	.v2c_parallelIn_1551(v2c_in1[155]),
	.v2c_parallelIn_1552(v2c_in2[155]),
	.v2c_parallelIn_1560(v2c_in0[156]),
	.v2c_parallelIn_1561(v2c_in1[156]),
	.v2c_parallelIn_1562(v2c_in2[156]),
	.v2c_parallelIn_1570(v2c_in0[157]),
	.v2c_parallelIn_1571(v2c_in1[157]),
	.v2c_parallelIn_1572(v2c_in2[157]),
	.v2c_parallelIn_1580(v2c_in0[158]),
	.v2c_parallelIn_1581(v2c_in1[158]),
	.v2c_parallelIn_1582(v2c_in2[158]),
	.v2c_parallelIn_1590(v2c_in0[159]),
	.v2c_parallelIn_1591(v2c_in1[159]),
	.v2c_parallelIn_1592(v2c_in2[159]),
	.v2c_parallelIn_1600(v2c_in0[160]),
	.v2c_parallelIn_1601(v2c_in1[160]),
	.v2c_parallelIn_1602(v2c_in2[160]),
	.v2c_parallelIn_1610(v2c_in0[161]),
	.v2c_parallelIn_1611(v2c_in1[161]),
	.v2c_parallelIn_1612(v2c_in2[161]),
	.v2c_parallelIn_1620(v2c_in0[162]),
	.v2c_parallelIn_1621(v2c_in1[162]),
	.v2c_parallelIn_1622(v2c_in2[162]),
	.v2c_parallelIn_1630(v2c_in0[163]),
	.v2c_parallelIn_1631(v2c_in1[163]),
	.v2c_parallelIn_1632(v2c_in2[163]),
	.v2c_parallelIn_1640(v2c_in0[164]),
	.v2c_parallelIn_1641(v2c_in1[164]),
	.v2c_parallelIn_1642(v2c_in2[164]),
	.v2c_parallelIn_1650(v2c_in0[165]),
	.v2c_parallelIn_1651(v2c_in1[165]),
	.v2c_parallelIn_1652(v2c_in2[165]),
	.v2c_parallelIn_1660(v2c_in0[166]),
	.v2c_parallelIn_1661(v2c_in1[166]),
	.v2c_parallelIn_1662(v2c_in2[166]),
	.v2c_parallelIn_1670(v2c_in0[167]),
	.v2c_parallelIn_1671(v2c_in1[167]),
	.v2c_parallelIn_1672(v2c_in2[167]),
	.v2c_parallelIn_1680(v2c_in0[168]),
	.v2c_parallelIn_1681(v2c_in1[168]),
	.v2c_parallelIn_1682(v2c_in2[168]),
	.v2c_parallelIn_1690(v2c_in0[169]),
	.v2c_parallelIn_1691(v2c_in1[169]),
	.v2c_parallelIn_1692(v2c_in2[169]),
	.v2c_parallelIn_1700(v2c_in0[170]),
	.v2c_parallelIn_1701(v2c_in1[170]),
	.v2c_parallelIn_1702(v2c_in2[170]),
	.v2c_parallelIn_1710(v2c_in0[171]),
	.v2c_parallelIn_1711(v2c_in1[171]),
	.v2c_parallelIn_1712(v2c_in2[171]),
	.v2c_parallelIn_1720(v2c_in0[172]),
	.v2c_parallelIn_1721(v2c_in1[172]),
	.v2c_parallelIn_1722(v2c_in2[172]),
	.v2c_parallelIn_1730(v2c_in0[173]),
	.v2c_parallelIn_1731(v2c_in1[173]),
	.v2c_parallelIn_1732(v2c_in2[173]),
	.v2c_parallelIn_1740(v2c_in0[174]),
	.v2c_parallelIn_1741(v2c_in1[174]),
	.v2c_parallelIn_1742(v2c_in2[174]),
	.v2c_parallelIn_1750(v2c_in0[175]),
	.v2c_parallelIn_1751(v2c_in1[175]),
	.v2c_parallelIn_1752(v2c_in2[175]),
	.v2c_parallelIn_1760(v2c_in0[176]),
	.v2c_parallelIn_1761(v2c_in1[176]),
	.v2c_parallelIn_1762(v2c_in2[176]),
	.v2c_parallelIn_1770(v2c_in0[177]),
	.v2c_parallelIn_1771(v2c_in1[177]),
	.v2c_parallelIn_1772(v2c_in2[177]),
	.v2c_parallelIn_1780(v2c_in0[178]),
	.v2c_parallelIn_1781(v2c_in1[178]),
	.v2c_parallelIn_1782(v2c_in2[178]),
	.v2c_parallelIn_1790(v2c_in0[179]),
	.v2c_parallelIn_1791(v2c_in1[179]),
	.v2c_parallelIn_1792(v2c_in2[179]),
	.v2c_parallelIn_1800(v2c_in0[180]),
	.v2c_parallelIn_1801(v2c_in1[180]),
	.v2c_parallelIn_1802(v2c_in2[180]),
	.v2c_parallelIn_1810(v2c_in0[181]),
	.v2c_parallelIn_1811(v2c_in1[181]),
	.v2c_parallelIn_1812(v2c_in2[181]),
	.v2c_parallelIn_1820(v2c_in0[182]),
	.v2c_parallelIn_1821(v2c_in1[182]),
	.v2c_parallelIn_1822(v2c_in2[182]),
	.v2c_parallelIn_1830(v2c_in0[183]),
	.v2c_parallelIn_1831(v2c_in1[183]),
	.v2c_parallelIn_1832(v2c_in2[183]),
	.v2c_parallelIn_1840(v2c_in0[184]),
	.v2c_parallelIn_1841(v2c_in1[184]),
	.v2c_parallelIn_1842(v2c_in2[184]),
	.v2c_parallelIn_1850(v2c_in0[185]),
	.v2c_parallelIn_1851(v2c_in1[185]),
	.v2c_parallelIn_1852(v2c_in2[185]),
	.v2c_parallelIn_1860(v2c_in0[186]),
	.v2c_parallelIn_1861(v2c_in1[186]),
	.v2c_parallelIn_1862(v2c_in2[186]),
	.v2c_parallelIn_1870(v2c_in0[187]),
	.v2c_parallelIn_1871(v2c_in1[187]),
	.v2c_parallelIn_1872(v2c_in2[187]),
	.v2c_parallelIn_1880(v2c_in0[188]),
	.v2c_parallelIn_1881(v2c_in1[188]),
	.v2c_parallelIn_1882(v2c_in2[188]),
	.v2c_parallelIn_1890(v2c_in0[189]),
	.v2c_parallelIn_1891(v2c_in1[189]),
	.v2c_parallelIn_1892(v2c_in2[189]),
	.v2c_parallelIn_1900(v2c_in0[190]),
	.v2c_parallelIn_1901(v2c_in1[190]),
	.v2c_parallelIn_1902(v2c_in2[190]),
	.v2c_parallelIn_1910(v2c_in0[191]),
	.v2c_parallelIn_1911(v2c_in1[191]),
	.v2c_parallelIn_1912(v2c_in2[191]),
	.v2c_parallelIn_1920(v2c_in0[192]),
	.v2c_parallelIn_1921(v2c_in1[192]),
	.v2c_parallelIn_1922(v2c_in2[192]),
	.v2c_parallelIn_1930(v2c_in0[193]),
	.v2c_parallelIn_1931(v2c_in1[193]),
	.v2c_parallelIn_1932(v2c_in2[193]),
	.v2c_parallelIn_1940(v2c_in0[194]),
	.v2c_parallelIn_1941(v2c_in1[194]),
	.v2c_parallelIn_1942(v2c_in2[194]),
	.v2c_parallelIn_1950(v2c_in0[195]),
	.v2c_parallelIn_1951(v2c_in1[195]),
	.v2c_parallelIn_1952(v2c_in2[195]),
	.v2c_parallelIn_1960(v2c_in0[196]),
	.v2c_parallelIn_1961(v2c_in1[196]),
	.v2c_parallelIn_1962(v2c_in2[196]),
	.v2c_parallelIn_1970(v2c_in0[197]),
	.v2c_parallelIn_1971(v2c_in1[197]),
	.v2c_parallelIn_1972(v2c_in2[197]),
	.v2c_parallelIn_1980(v2c_in0[198]),
	.v2c_parallelIn_1981(v2c_in1[198]),
	.v2c_parallelIn_1982(v2c_in2[198]),
	.v2c_parallelIn_1990(v2c_in0[199]),
	.v2c_parallelIn_1991(v2c_in1[199]),
	.v2c_parallelIn_1992(v2c_in2[199]),
	.v2c_parallelIn_2000(v2c_in0[200]),
	.v2c_parallelIn_2001(v2c_in1[200]),
	.v2c_parallelIn_2002(v2c_in2[200]),
	.v2c_parallelIn_2010(v2c_in0[201]),
	.v2c_parallelIn_2011(v2c_in1[201]),
	.v2c_parallelIn_2012(v2c_in2[201]),
	.v2c_parallelIn_2020(v2c_in0[202]),
	.v2c_parallelIn_2021(v2c_in1[202]),
	.v2c_parallelIn_2022(v2c_in2[202]),
	.v2c_parallelIn_2030(v2c_in0[203]),
	.v2c_parallelIn_2031(v2c_in1[203]),
	.v2c_parallelIn_2032(v2c_in2[203]),
	
	.load(load[1:0]),
	.parallel_en (parallel_en[1:0]),
	.serial_clk (read_clk)
);
endmodule