module qsn_merge (
	output wire [254:0] sw_out,

	input wire [253:0] left_in,
	input wire [254:0] right_in,
	input wire [253:0] sel
);

	assign sw_out[0] = (sel[0] == 1'b0) ? right_in[254] : left_in[0];
	assign sw_out[1] = (sel[1] == 1'b0) ? right_in[253] : left_in[1];
	assign sw_out[2] = (sel[2] == 1'b0) ? right_in[252] : left_in[2];
	assign sw_out[3] = (sel[3] == 1'b0) ? right_in[251] : left_in[3];
	assign sw_out[4] = (sel[4] == 1'b0) ? right_in[250] : left_in[4];
	assign sw_out[5] = (sel[5] == 1'b0) ? right_in[249] : left_in[5];
	assign sw_out[6] = (sel[6] == 1'b0) ? right_in[248] : left_in[6];
	assign sw_out[7] = (sel[7] == 1'b0) ? right_in[247] : left_in[7];
	assign sw_out[8] = (sel[8] == 1'b0) ? right_in[246] : left_in[8];
	assign sw_out[9] = (sel[9] == 1'b0) ? right_in[245] : left_in[9];
	assign sw_out[10] = (sel[10] == 1'b0) ? right_in[244] : left_in[10];
	assign sw_out[11] = (sel[11] == 1'b0) ? right_in[243] : left_in[11];
	assign sw_out[12] = (sel[12] == 1'b0) ? right_in[242] : left_in[12];
	assign sw_out[13] = (sel[13] == 1'b0) ? right_in[241] : left_in[13];
	assign sw_out[14] = (sel[14] == 1'b0) ? right_in[240] : left_in[14];
	assign sw_out[15] = (sel[15] == 1'b0) ? right_in[239] : left_in[15];
	assign sw_out[16] = (sel[16] == 1'b0) ? right_in[238] : left_in[16];
	assign sw_out[17] = (sel[17] == 1'b0) ? right_in[237] : left_in[17];
	assign sw_out[18] = (sel[18] == 1'b0) ? right_in[236] : left_in[18];
	assign sw_out[19] = (sel[19] == 1'b0) ? right_in[235] : left_in[19];
	assign sw_out[20] = (sel[20] == 1'b0) ? right_in[234] : left_in[20];
	assign sw_out[21] = (sel[21] == 1'b0) ? right_in[233] : left_in[21];
	assign sw_out[22] = (sel[22] == 1'b0) ? right_in[232] : left_in[22];
	assign sw_out[23] = (sel[23] == 1'b0) ? right_in[231] : left_in[23];
	assign sw_out[24] = (sel[24] == 1'b0) ? right_in[230] : left_in[24];
	assign sw_out[25] = (sel[25] == 1'b0) ? right_in[229] : left_in[25];
	assign sw_out[26] = (sel[26] == 1'b0) ? right_in[228] : left_in[26];
	assign sw_out[27] = (sel[27] == 1'b0) ? right_in[227] : left_in[27];
	assign sw_out[28] = (sel[28] == 1'b0) ? right_in[226] : left_in[28];
	assign sw_out[29] = (sel[29] == 1'b0) ? right_in[225] : left_in[29];
	assign sw_out[30] = (sel[30] == 1'b0) ? right_in[224] : left_in[30];
	assign sw_out[31] = (sel[31] == 1'b0) ? right_in[223] : left_in[31];
	assign sw_out[32] = (sel[32] == 1'b0) ? right_in[222] : left_in[32];
	assign sw_out[33] = (sel[33] == 1'b0) ? right_in[221] : left_in[33];
	assign sw_out[34] = (sel[34] == 1'b0) ? right_in[220] : left_in[34];
	assign sw_out[35] = (sel[35] == 1'b0) ? right_in[219] : left_in[35];
	assign sw_out[36] = (sel[36] == 1'b0) ? right_in[218] : left_in[36];
	assign sw_out[37] = (sel[37] == 1'b0) ? right_in[217] : left_in[37];
	assign sw_out[38] = (sel[38] == 1'b0) ? right_in[216] : left_in[38];
	assign sw_out[39] = (sel[39] == 1'b0) ? right_in[215] : left_in[39];
	assign sw_out[40] = (sel[40] == 1'b0) ? right_in[214] : left_in[40];
	assign sw_out[41] = (sel[41] == 1'b0) ? right_in[213] : left_in[41];
	assign sw_out[42] = (sel[42] == 1'b0) ? right_in[212] : left_in[42];
	assign sw_out[43] = (sel[43] == 1'b0) ? right_in[211] : left_in[43];
	assign sw_out[44] = (sel[44] == 1'b0) ? right_in[210] : left_in[44];
	assign sw_out[45] = (sel[45] == 1'b0) ? right_in[209] : left_in[45];
	assign sw_out[46] = (sel[46] == 1'b0) ? right_in[208] : left_in[46];
	assign sw_out[47] = (sel[47] == 1'b0) ? right_in[207] : left_in[47];
	assign sw_out[48] = (sel[48] == 1'b0) ? right_in[206] : left_in[48];
	assign sw_out[49] = (sel[49] == 1'b0) ? right_in[205] : left_in[49];
	assign sw_out[50] = (sel[50] == 1'b0) ? right_in[204] : left_in[50];
	assign sw_out[51] = (sel[51] == 1'b0) ? right_in[203] : left_in[51];
	assign sw_out[52] = (sel[52] == 1'b0) ? right_in[202] : left_in[52];
	assign sw_out[53] = (sel[53] == 1'b0) ? right_in[201] : left_in[53];
	assign sw_out[54] = (sel[54] == 1'b0) ? right_in[200] : left_in[54];
	assign sw_out[55] = (sel[55] == 1'b0) ? right_in[199] : left_in[55];
	assign sw_out[56] = (sel[56] == 1'b0) ? right_in[198] : left_in[56];
	assign sw_out[57] = (sel[57] == 1'b0) ? right_in[197] : left_in[57];
	assign sw_out[58] = (sel[58] == 1'b0) ? right_in[196] : left_in[58];
	assign sw_out[59] = (sel[59] == 1'b0) ? right_in[195] : left_in[59];
	assign sw_out[60] = (sel[60] == 1'b0) ? right_in[194] : left_in[60];
	assign sw_out[61] = (sel[61] == 1'b0) ? right_in[193] : left_in[61];
	assign sw_out[62] = (sel[62] == 1'b0) ? right_in[192] : left_in[62];
	assign sw_out[63] = (sel[63] == 1'b0) ? right_in[191] : left_in[63];
	assign sw_out[64] = (sel[64] == 1'b0) ? right_in[190] : left_in[64];
	assign sw_out[65] = (sel[65] == 1'b0) ? right_in[189] : left_in[65];
	assign sw_out[66] = (sel[66] == 1'b0) ? right_in[188] : left_in[66];
	assign sw_out[67] = (sel[67] == 1'b0) ? right_in[187] : left_in[67];
	assign sw_out[68] = (sel[68] == 1'b0) ? right_in[186] : left_in[68];
	assign sw_out[69] = (sel[69] == 1'b0) ? right_in[185] : left_in[69];
	assign sw_out[70] = (sel[70] == 1'b0) ? right_in[184] : left_in[70];
	assign sw_out[71] = (sel[71] == 1'b0) ? right_in[183] : left_in[71];
	assign sw_out[72] = (sel[72] == 1'b0) ? right_in[182] : left_in[72];
	assign sw_out[73] = (sel[73] == 1'b0) ? right_in[181] : left_in[73];
	assign sw_out[74] = (sel[74] == 1'b0) ? right_in[180] : left_in[74];
	assign sw_out[75] = (sel[75] == 1'b0) ? right_in[179] : left_in[75];
	assign sw_out[76] = (sel[76] == 1'b0) ? right_in[178] : left_in[76];
	assign sw_out[77] = (sel[77] == 1'b0) ? right_in[177] : left_in[77];
	assign sw_out[78] = (sel[78] == 1'b0) ? right_in[176] : left_in[78];
	assign sw_out[79] = (sel[79] == 1'b0) ? right_in[175] : left_in[79];
	assign sw_out[80] = (sel[80] == 1'b0) ? right_in[174] : left_in[80];
	assign sw_out[81] = (sel[81] == 1'b0) ? right_in[173] : left_in[81];
	assign sw_out[82] = (sel[82] == 1'b0) ? right_in[172] : left_in[82];
	assign sw_out[83] = (sel[83] == 1'b0) ? right_in[171] : left_in[83];
	assign sw_out[84] = (sel[84] == 1'b0) ? right_in[170] : left_in[84];
	assign sw_out[85] = (sel[85] == 1'b0) ? right_in[169] : left_in[85];
	assign sw_out[86] = (sel[86] == 1'b0) ? right_in[168] : left_in[86];
	assign sw_out[87] = (sel[87] == 1'b0) ? right_in[167] : left_in[87];
	assign sw_out[88] = (sel[88] == 1'b0) ? right_in[166] : left_in[88];
	assign sw_out[89] = (sel[89] == 1'b0) ? right_in[165] : left_in[89];
	assign sw_out[90] = (sel[90] == 1'b0) ? right_in[164] : left_in[90];
	assign sw_out[91] = (sel[91] == 1'b0) ? right_in[163] : left_in[91];
	assign sw_out[92] = (sel[92] == 1'b0) ? right_in[162] : left_in[92];
	assign sw_out[93] = (sel[93] == 1'b0) ? right_in[161] : left_in[93];
	assign sw_out[94] = (sel[94] == 1'b0) ? right_in[160] : left_in[94];
	assign sw_out[95] = (sel[95] == 1'b0) ? right_in[159] : left_in[95];
	assign sw_out[96] = (sel[96] == 1'b0) ? right_in[158] : left_in[96];
	assign sw_out[97] = (sel[97] == 1'b0) ? right_in[157] : left_in[97];
	assign sw_out[98] = (sel[98] == 1'b0) ? right_in[156] : left_in[98];
	assign sw_out[99] = (sel[99] == 1'b0) ? right_in[155] : left_in[99];
	assign sw_out[100] = (sel[100] == 1'b0) ? right_in[154] : left_in[100];
	assign sw_out[101] = (sel[101] == 1'b0) ? right_in[153] : left_in[101];
	assign sw_out[102] = (sel[102] == 1'b0) ? right_in[152] : left_in[102];
	assign sw_out[103] = (sel[103] == 1'b0) ? right_in[151] : left_in[103];
	assign sw_out[104] = (sel[104] == 1'b0) ? right_in[150] : left_in[104];
	assign sw_out[105] = (sel[105] == 1'b0) ? right_in[149] : left_in[105];
	assign sw_out[106] = (sel[106] == 1'b0) ? right_in[148] : left_in[106];
	assign sw_out[107] = (sel[107] == 1'b0) ? right_in[147] : left_in[107];
	assign sw_out[108] = (sel[108] == 1'b0) ? right_in[146] : left_in[108];
	assign sw_out[109] = (sel[109] == 1'b0) ? right_in[145] : left_in[109];
	assign sw_out[110] = (sel[110] == 1'b0) ? right_in[144] : left_in[110];
	assign sw_out[111] = (sel[111] == 1'b0) ? right_in[143] : left_in[111];
	assign sw_out[112] = (sel[112] == 1'b0) ? right_in[142] : left_in[112];
	assign sw_out[113] = (sel[113] == 1'b0) ? right_in[141] : left_in[113];
	assign sw_out[114] = (sel[114] == 1'b0) ? right_in[140] : left_in[114];
	assign sw_out[115] = (sel[115] == 1'b0) ? right_in[139] : left_in[115];
	assign sw_out[116] = (sel[116] == 1'b0) ? right_in[138] : left_in[116];
	assign sw_out[117] = (sel[117] == 1'b0) ? right_in[137] : left_in[117];
	assign sw_out[118] = (sel[118] == 1'b0) ? right_in[136] : left_in[118];
	assign sw_out[119] = (sel[119] == 1'b0) ? right_in[135] : left_in[119];
	assign sw_out[120] = (sel[120] == 1'b0) ? right_in[134] : left_in[120];
	assign sw_out[121] = (sel[121] == 1'b0) ? right_in[133] : left_in[121];
	assign sw_out[122] = (sel[122] == 1'b0) ? right_in[132] : left_in[122];
	assign sw_out[123] = (sel[123] == 1'b0) ? right_in[131] : left_in[123];
	assign sw_out[124] = (sel[124] == 1'b0) ? right_in[130] : left_in[124];
	assign sw_out[125] = (sel[125] == 1'b0) ? right_in[129] : left_in[125];
	assign sw_out[126] = (sel[126] == 1'b0) ? right_in[128] : left_in[126];
	assign sw_out[127] = (sel[127] == 1'b0) ? right_in[127] : left_in[127];
	assign sw_out[128] = (sel[128] == 1'b0) ? right_in[126] : left_in[128];
	assign sw_out[129] = (sel[129] == 1'b0) ? right_in[125] : left_in[129];
	assign sw_out[130] = (sel[130] == 1'b0) ? right_in[124] : left_in[130];
	assign sw_out[131] = (sel[131] == 1'b0) ? right_in[123] : left_in[131];
	assign sw_out[132] = (sel[132] == 1'b0) ? right_in[122] : left_in[132];
	assign sw_out[133] = (sel[133] == 1'b0) ? right_in[121] : left_in[133];
	assign sw_out[134] = (sel[134] == 1'b0) ? right_in[120] : left_in[134];
	assign sw_out[135] = (sel[135] == 1'b0) ? right_in[119] : left_in[135];
	assign sw_out[136] = (sel[136] == 1'b0) ? right_in[118] : left_in[136];
	assign sw_out[137] = (sel[137] == 1'b0) ? right_in[117] : left_in[137];
	assign sw_out[138] = (sel[138] == 1'b0) ? right_in[116] : left_in[138];
	assign sw_out[139] = (sel[139] == 1'b0) ? right_in[115] : left_in[139];
	assign sw_out[140] = (sel[140] == 1'b0) ? right_in[114] : left_in[140];
	assign sw_out[141] = (sel[141] == 1'b0) ? right_in[113] : left_in[141];
	assign sw_out[142] = (sel[142] == 1'b0) ? right_in[112] : left_in[142];
	assign sw_out[143] = (sel[143] == 1'b0) ? right_in[111] : left_in[143];
	assign sw_out[144] = (sel[144] == 1'b0) ? right_in[110] : left_in[144];
	assign sw_out[145] = (sel[145] == 1'b0) ? right_in[109] : left_in[145];
	assign sw_out[146] = (sel[146] == 1'b0) ? right_in[108] : left_in[146];
	assign sw_out[147] = (sel[147] == 1'b0) ? right_in[107] : left_in[147];
	assign sw_out[148] = (sel[148] == 1'b0) ? right_in[106] : left_in[148];
	assign sw_out[149] = (sel[149] == 1'b0) ? right_in[105] : left_in[149];
	assign sw_out[150] = (sel[150] == 1'b0) ? right_in[104] : left_in[150];
	assign sw_out[151] = (sel[151] == 1'b0) ? right_in[103] : left_in[151];
	assign sw_out[152] = (sel[152] == 1'b0) ? right_in[102] : left_in[152];
	assign sw_out[153] = (sel[153] == 1'b0) ? right_in[101] : left_in[153];
	assign sw_out[154] = (sel[154] == 1'b0) ? right_in[100] : left_in[154];
	assign sw_out[155] = (sel[155] == 1'b0) ? right_in[99] : left_in[155];
	assign sw_out[156] = (sel[156] == 1'b0) ? right_in[98] : left_in[156];
	assign sw_out[157] = (sel[157] == 1'b0) ? right_in[97] : left_in[157];
	assign sw_out[158] = (sel[158] == 1'b0) ? right_in[96] : left_in[158];
	assign sw_out[159] = (sel[159] == 1'b0) ? right_in[95] : left_in[159];
	assign sw_out[160] = (sel[160] == 1'b0) ? right_in[94] : left_in[160];
	assign sw_out[161] = (sel[161] == 1'b0) ? right_in[93] : left_in[161];
	assign sw_out[162] = (sel[162] == 1'b0) ? right_in[92] : left_in[162];
	assign sw_out[163] = (sel[163] == 1'b0) ? right_in[91] : left_in[163];
	assign sw_out[164] = (sel[164] == 1'b0) ? right_in[90] : left_in[164];
	assign sw_out[165] = (sel[165] == 1'b0) ? right_in[89] : left_in[165];
	assign sw_out[166] = (sel[166] == 1'b0) ? right_in[88] : left_in[166];
	assign sw_out[167] = (sel[167] == 1'b0) ? right_in[87] : left_in[167];
	assign sw_out[168] = (sel[168] == 1'b0) ? right_in[86] : left_in[168];
	assign sw_out[169] = (sel[169] == 1'b0) ? right_in[85] : left_in[169];
	assign sw_out[170] = (sel[170] == 1'b0) ? right_in[84] : left_in[170];
	assign sw_out[171] = (sel[171] == 1'b0) ? right_in[83] : left_in[171];
	assign sw_out[172] = (sel[172] == 1'b0) ? right_in[82] : left_in[172];
	assign sw_out[173] = (sel[173] == 1'b0) ? right_in[81] : left_in[173];
	assign sw_out[174] = (sel[174] == 1'b0) ? right_in[80] : left_in[174];
	assign sw_out[175] = (sel[175] == 1'b0) ? right_in[79] : left_in[175];
	assign sw_out[176] = (sel[176] == 1'b0) ? right_in[78] : left_in[176];
	assign sw_out[177] = (sel[177] == 1'b0) ? right_in[77] : left_in[177];
	assign sw_out[178] = (sel[178] == 1'b0) ? right_in[76] : left_in[178];
	assign sw_out[179] = (sel[179] == 1'b0) ? right_in[75] : left_in[179];
	assign sw_out[180] = (sel[180] == 1'b0) ? right_in[74] : left_in[180];
	assign sw_out[181] = (sel[181] == 1'b0) ? right_in[73] : left_in[181];
	assign sw_out[182] = (sel[182] == 1'b0) ? right_in[72] : left_in[182];
	assign sw_out[183] = (sel[183] == 1'b0) ? right_in[71] : left_in[183];
	assign sw_out[184] = (sel[184] == 1'b0) ? right_in[70] : left_in[184];
	assign sw_out[185] = (sel[185] == 1'b0) ? right_in[69] : left_in[185];
	assign sw_out[186] = (sel[186] == 1'b0) ? right_in[68] : left_in[186];
	assign sw_out[187] = (sel[187] == 1'b0) ? right_in[67] : left_in[187];
	assign sw_out[188] = (sel[188] == 1'b0) ? right_in[66] : left_in[188];
	assign sw_out[189] = (sel[189] == 1'b0) ? right_in[65] : left_in[189];
	assign sw_out[190] = (sel[190] == 1'b0) ? right_in[64] : left_in[190];
	assign sw_out[191] = (sel[191] == 1'b0) ? right_in[63] : left_in[191];
	assign sw_out[192] = (sel[192] == 1'b0) ? right_in[62] : left_in[192];
	assign sw_out[193] = (sel[193] == 1'b0) ? right_in[61] : left_in[193];
	assign sw_out[194] = (sel[194] == 1'b0) ? right_in[60] : left_in[194];
	assign sw_out[195] = (sel[195] == 1'b0) ? right_in[59] : left_in[195];
	assign sw_out[196] = (sel[196] == 1'b0) ? right_in[58] : left_in[196];
	assign sw_out[197] = (sel[197] == 1'b0) ? right_in[57] : left_in[197];
	assign sw_out[198] = (sel[198] == 1'b0) ? right_in[56] : left_in[198];
	assign sw_out[199] = (sel[199] == 1'b0) ? right_in[55] : left_in[199];
	assign sw_out[200] = (sel[200] == 1'b0) ? right_in[54] : left_in[200];
	assign sw_out[201] = (sel[201] == 1'b0) ? right_in[53] : left_in[201];
	assign sw_out[202] = (sel[202] == 1'b0) ? right_in[52] : left_in[202];
	assign sw_out[203] = (sel[203] == 1'b0) ? right_in[51] : left_in[203];
	assign sw_out[204] = (sel[204] == 1'b0) ? right_in[50] : left_in[204];
	assign sw_out[205] = (sel[205] == 1'b0) ? right_in[49] : left_in[205];
	assign sw_out[206] = (sel[206] == 1'b0) ? right_in[48] : left_in[206];
	assign sw_out[207] = (sel[207] == 1'b0) ? right_in[47] : left_in[207];
	assign sw_out[208] = (sel[208] == 1'b0) ? right_in[46] : left_in[208];
	assign sw_out[209] = (sel[209] == 1'b0) ? right_in[45] : left_in[209];
	assign sw_out[210] = (sel[210] == 1'b0) ? right_in[44] : left_in[210];
	assign sw_out[211] = (sel[211] == 1'b0) ? right_in[43] : left_in[211];
	assign sw_out[212] = (sel[212] == 1'b0) ? right_in[42] : left_in[212];
	assign sw_out[213] = (sel[213] == 1'b0) ? right_in[41] : left_in[213];
	assign sw_out[214] = (sel[214] == 1'b0) ? right_in[40] : left_in[214];
	assign sw_out[215] = (sel[215] == 1'b0) ? right_in[39] : left_in[215];
	assign sw_out[216] = (sel[216] == 1'b0) ? right_in[38] : left_in[216];
	assign sw_out[217] = (sel[217] == 1'b0) ? right_in[37] : left_in[217];
	assign sw_out[218] = (sel[218] == 1'b0) ? right_in[36] : left_in[218];
	assign sw_out[219] = (sel[219] == 1'b0) ? right_in[35] : left_in[219];
	assign sw_out[220] = (sel[220] == 1'b0) ? right_in[34] : left_in[220];
	assign sw_out[221] = (sel[221] == 1'b0) ? right_in[33] : left_in[221];
	assign sw_out[222] = (sel[222] == 1'b0) ? right_in[32] : left_in[222];
	assign sw_out[223] = (sel[223] == 1'b0) ? right_in[31] : left_in[223];
	assign sw_out[224] = (sel[224] == 1'b0) ? right_in[30] : left_in[224];
	assign sw_out[225] = (sel[225] == 1'b0) ? right_in[29] : left_in[225];
	assign sw_out[226] = (sel[226] == 1'b0) ? right_in[28] : left_in[226];
	assign sw_out[227] = (sel[227] == 1'b0) ? right_in[27] : left_in[227];
	assign sw_out[228] = (sel[228] == 1'b0) ? right_in[26] : left_in[228];
	assign sw_out[229] = (sel[229] == 1'b0) ? right_in[25] : left_in[229];
	assign sw_out[230] = (sel[230] == 1'b0) ? right_in[24] : left_in[230];
	assign sw_out[231] = (sel[231] == 1'b0) ? right_in[23] : left_in[231];
	assign sw_out[232] = (sel[232] == 1'b0) ? right_in[22] : left_in[232];
	assign sw_out[233] = (sel[233] == 1'b0) ? right_in[21] : left_in[233];
	assign sw_out[234] = (sel[234] == 1'b0) ? right_in[20] : left_in[234];
	assign sw_out[235] = (sel[235] == 1'b0) ? right_in[19] : left_in[235];
	assign sw_out[236] = (sel[236] == 1'b0) ? right_in[18] : left_in[236];
	assign sw_out[237] = (sel[237] == 1'b0) ? right_in[17] : left_in[237];
	assign sw_out[238] = (sel[238] == 1'b0) ? right_in[16] : left_in[238];
	assign sw_out[239] = (sel[239] == 1'b0) ? right_in[15] : left_in[239];
	assign sw_out[240] = (sel[240] == 1'b0) ? right_in[14] : left_in[240];
	assign sw_out[241] = (sel[241] == 1'b0) ? right_in[13] : left_in[241];
	assign sw_out[242] = (sel[242] == 1'b0) ? right_in[12] : left_in[242];
	assign sw_out[243] = (sel[243] == 1'b0) ? right_in[11] : left_in[243];
	assign sw_out[244] = (sel[244] == 1'b0) ? right_in[10] : left_in[244];
	assign sw_out[245] = (sel[245] == 1'b0) ? right_in[9] : left_in[245];
	assign sw_out[246] = (sel[246] == 1'b0) ? right_in[8] : left_in[246];
	assign sw_out[247] = (sel[247] == 1'b0) ? right_in[7] : left_in[247];
	assign sw_out[248] = (sel[248] == 1'b0) ? right_in[6] : left_in[248];
	assign sw_out[249] = (sel[249] == 1'b0) ? right_in[5] : left_in[249];
	assign sw_out[250] = (sel[250] == 1'b0) ? right_in[4] : left_in[250];
	assign sw_out[251] = (sel[251] == 1'b0) ? right_in[3] : left_in[251];
	assign sw_out[252] = (sel[252] == 1'b0) ? right_in[2] : left_in[252];
	assign sw_out[253] = (sel[253] == 1'b0) ? right_in[1] : left_in[253];
	assign sw_out[254] = right_in[0];
endmodule