module test #(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 85,
	parameter RAM_UNIT_MSG_NUM = 17, // each RAM unit contributes 17 messages of size 4-bit
	parameter RAM_PORTA_RANGE = 9, // 9 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port A,
	parameter RAM_PORTB_RANGE = 8, // 8 out of RAM_UNIT_MSG_NUM messages are from/to true dual-port of RAM unit port b, 
	parameter MEM_DEVICE_NUM = 5,
	parameter DEPTH = 1024,
	parameter WIDTH = 36,
	parameter ADDR = $clog2(DEPTH)
)(
	output wire Dout,

	input wire [QUAN_SIZE-1:0] Din,
	input wire [ADDR-1:0] sync_addr,
	input wire we,
	input wire sys_clk
);

wire [QUAN_SIZE-1:0] dout_reg [0:CHECK_PARALLELISM-1];
	column_ram_pc85 #(
			.QUAN_SIZE(QUAN_SIZE),
			.CHECK_PARALLELISM(CHECK_PARALLELISM),
			.RAM_UNIT_MSG_NUM(RAM_UNIT_MSG_NUM),
			.RAM_PORTA_RANGE(RAM_PORTA_RANGE),
			.RAM_PORTB_RANGE(RAM_PORTB_RANGE),
			.MEM_DEVICE_NUM(MEM_DEVICE_NUM),
			.DEPTH(DEPTH),
			.WIDTH(WIDTH),
			.ADDR(ADDR)
		) inst_column_ram_pc85 (
		.Dout_0	(dout_reg[0]),
		.Dout_1	(dout_reg[1]),
		.Dout_2	(dout_reg[2]),
		.Dout_3	(dout_reg[3]),
		.Dout_4	(dout_reg[4]),
		.Dout_5	(dout_reg[5]),
		.Dout_6	(dout_reg[6]),
		.Dout_7	(dout_reg[7]),
		.Dout_8	(dout_reg[8]),
		.Dout_9	(dout_reg[9]),
		.Dout_10	(dout_reg[10]),
		.Dout_11	(dout_reg[11]),
		.Dout_12	(dout_reg[12]),
		.Dout_13	(dout_reg[13]),
		.Dout_14	(dout_reg[14]),
		.Dout_15	(dout_reg[15]),
		.Dout_16	(dout_reg[16]),
		.Dout_17	(dout_reg[17]),
		.Dout_18	(dout_reg[18]),
		.Dout_19	(dout_reg[19]),
		.Dout_20	(dout_reg[20]),
		.Dout_21	(dout_reg[21]),
		.Dout_22	(dout_reg[22]),
		.Dout_23	(dout_reg[23]),
		.Dout_24	(dout_reg[24]),
		.Dout_25	(dout_reg[25]),
		.Dout_26	(dout_reg[26]),
		.Dout_27	(dout_reg[27]),
		.Dout_28	(dout_reg[28]),
		.Dout_29	(dout_reg[29]),
		.Dout_30	(dout_reg[30]),
		.Dout_31	(dout_reg[31]),
		.Dout_32	(dout_reg[32]),
		.Dout_33	(dout_reg[33]),
		.Dout_34	(dout_reg[34]),
		.Dout_35	(dout_reg[35]),
		.Dout_36	(dout_reg[36]),
		.Dout_37	(dout_reg[37]),
		.Dout_38	(dout_reg[38]),
		.Dout_39	(dout_reg[39]),
		.Dout_40	(dout_reg[40]),
		.Dout_41	(dout_reg[41]),
		.Dout_42	(dout_reg[42]),
		.Dout_43	(dout_reg[43]),
		.Dout_44	(dout_reg[44]),
		.Dout_45	(dout_reg[45]),
		.Dout_46	(dout_reg[46]),
		.Dout_47	(dout_reg[47]),
		.Dout_48	(dout_reg[48]),
		.Dout_49	(dout_reg[49]),
		.Dout_50	(dout_reg[50]),
		.Dout_51	(dout_reg[51]),
		.Dout_52	(dout_reg[52]),
		.Dout_53	(dout_reg[53]),
		.Dout_54	(dout_reg[54]),
		.Dout_55	(dout_reg[55]),
		.Dout_56	(dout_reg[56]),
		.Dout_57	(dout_reg[57]),
		.Dout_58	(dout_reg[58]),
		.Dout_59	(dout_reg[59]),
		.Dout_60	(dout_reg[60]),
		.Dout_61	(dout_reg[61]),
		.Dout_62	(dout_reg[62]),
		.Dout_63	(dout_reg[63]),
		.Dout_64	(dout_reg[64]),
		.Dout_65	(dout_reg[65]),
		.Dout_66	(dout_reg[66]),
		.Dout_67	(dout_reg[67]),
		.Dout_68	(dout_reg[68]),
		.Dout_69	(dout_reg[69]),
		.Dout_70	(dout_reg[70]),
		.Dout_71	(dout_reg[71]),
		.Dout_72	(dout_reg[72]),
		.Dout_73	(dout_reg[73]),
		.Dout_74	(dout_reg[74]),
		.Dout_75	(dout_reg[75]),
		.Dout_76	(dout_reg[76]),
		.Dout_77	(dout_reg[77]),
		.Dout_78	(dout_reg[78]),
		.Dout_79	(dout_reg[79]),
		.Dout_80	(dout_reg[80]),
		.Dout_81	(dout_reg[81]),
		.Dout_82	(dout_reg[82]),
		.Dout_83	(dout_reg[83]),
		.Dout_84	(dout_reg[84]),

			.Din_0     (Din[QUAN_SIZE-1:0]),
			.Din_1     (Din[QUAN_SIZE-1:0]),
			.Din_2     (Din[QUAN_SIZE-1:0]),
			.Din_3     (Din[QUAN_SIZE-1:0]),
			.Din_4     (Din[QUAN_SIZE-1:0]),
			.Din_5     (Din[QUAN_SIZE-1:0]),
			.Din_6     (Din[QUAN_SIZE-1:0]),
			.Din_7     (Din[QUAN_SIZE-1:0]),
			.Din_8     (Din[QUAN_SIZE-1:0]),
			.Din_9     (Din[QUAN_SIZE-1:0]),
			.Din_10    (Din[QUAN_SIZE-1:0]),
			.Din_11    (Din[QUAN_SIZE-1:0]),
			.Din_12    (Din[QUAN_SIZE-1:0]),
			.Din_13    (Din[QUAN_SIZE-1:0]),
			.Din_14    (Din[QUAN_SIZE-1:0]),
			.Din_15    (Din[QUAN_SIZE-1:0]),
			.Din_16    (Din[QUAN_SIZE-1:0]),
			.Din_17    (Din[QUAN_SIZE-1:0]),
			.Din_18    (Din[QUAN_SIZE-1:0]),
			.Din_19    (Din[QUAN_SIZE-1:0]),
			.Din_20    (Din[QUAN_SIZE-1:0]),
			.Din_21    (Din[QUAN_SIZE-1:0]),
			.Din_22    (Din[QUAN_SIZE-1:0]),
			.Din_23    (Din[QUAN_SIZE-1:0]),
			.Din_24    (Din[QUAN_SIZE-1:0]),
			.Din_25    (Din[QUAN_SIZE-1:0]),
			.Din_26    (Din[QUAN_SIZE-1:0]),
			.Din_27    (Din[QUAN_SIZE-1:0]),
			.Din_28    (Din[QUAN_SIZE-1:0]),
			.Din_29    (Din[QUAN_SIZE-1:0]),
			.Din_30    (Din[QUAN_SIZE-1:0]),
			.Din_31    (Din[QUAN_SIZE-1:0]),
			.Din_32    (Din[QUAN_SIZE-1:0]),
			.Din_33    (Din[QUAN_SIZE-1:0]),
			.Din_34    (Din[QUAN_SIZE-1:0]),
			.Din_35    (Din[QUAN_SIZE-1:0]),
			.Din_36    (Din[QUAN_SIZE-1:0]),
			.Din_37    (Din[QUAN_SIZE-1:0]),
			.Din_38    (Din[QUAN_SIZE-1:0]),
			.Din_39    (Din[QUAN_SIZE-1:0]),
			.Din_40    (Din[QUAN_SIZE-1:0]),
			.Din_41    (Din[QUAN_SIZE-1:0]),
			.Din_42    (Din[QUAN_SIZE-1:0]),
			.Din_43    (Din[QUAN_SIZE-1:0]),
			.Din_44    (Din[QUAN_SIZE-1:0]),
			.Din_45    (Din[QUAN_SIZE-1:0]),
			.Din_46    (Din[QUAN_SIZE-1:0]),
			.Din_47    (Din[QUAN_SIZE-1:0]),
			.Din_48    (Din[QUAN_SIZE-1:0]),
			.Din_49    (Din[QUAN_SIZE-1:0]),
			.Din_50    (Din[QUAN_SIZE-1:0]),
			.Din_51    (Din[QUAN_SIZE-1:0]),
			.Din_52    (Din[QUAN_SIZE-1:0]),
			.Din_53    (Din[QUAN_SIZE-1:0]),
			.Din_54    (Din[QUAN_SIZE-1:0]),
			.Din_55    (Din[QUAN_SIZE-1:0]),
			.Din_56    (Din[QUAN_SIZE-1:0]),
			.Din_57    (Din[QUAN_SIZE-1:0]),
			.Din_58    (Din[QUAN_SIZE-1:0]),
			.Din_59    (Din[QUAN_SIZE-1:0]),
			.Din_60    (Din[QUAN_SIZE-1:0]),
			.Din_61    (Din[QUAN_SIZE-1:0]),
			.Din_62    (Din[QUAN_SIZE-1:0]),
			.Din_63    (Din[QUAN_SIZE-1:0]),
			.Din_64    (Din[QUAN_SIZE-1:0]),
			.Din_65    (Din[QUAN_SIZE-1:0]),
			.Din_66    (Din[QUAN_SIZE-1:0]),
			.Din_67    (Din[QUAN_SIZE-1:0]),
			.Din_68    (Din[QUAN_SIZE-1:0]),
			.Din_69    (Din[QUAN_SIZE-1:0]),
			.Din_70    (Din[QUAN_SIZE-1:0]),
			.Din_71    (Din[QUAN_SIZE-1:0]),
			.Din_72    (Din[QUAN_SIZE-1:0]),
			.Din_73    (Din[QUAN_SIZE-1:0]),
			.Din_74    (Din[QUAN_SIZE-1:0]),
			.Din_75    (Din[QUAN_SIZE-1:0]),
			.Din_76    (Din[QUAN_SIZE-1:0]),
			.Din_77    (Din[QUAN_SIZE-1:0]),
			.Din_78    (Din[QUAN_SIZE-1:0]),
			.Din_79    (Din[QUAN_SIZE-1:0]),
			.Din_80    (Din[QUAN_SIZE-1:0]),
			.Din_81    (Din[QUAN_SIZE-1:0]),
			.Din_82    (Din[QUAN_SIZE-1:0]),
			.Din_83    (Din[QUAN_SIZE-1:0]),
			.Din_84    (Din[QUAN_SIZE-1:0]),
			.sync_addr (sync_addr),
			.we        (we),
			.sys_clk   (sys_clk)
		);

	reductin_or reductin_or_u0 (
		.dout (Dout),
		.din_0 (dout_reg[0]),
		.din_1 (dout_reg[1]),
		.din_2 (dout_reg[2]),
		.din_3 (dout_reg[3]),
		.din_4 (dout_reg[4]),
		.din_5 (dout_reg[5]),
		.din_6 (dout_reg[6]),
		.din_7 (dout_reg[7]),
		.din_8 (dout_reg[8]),
		.din_9 (dout_reg[9]),
		.din_10 (dout_reg[10]),
		.din_11 (dout_reg[11]),
		.din_12 (dout_reg[12]),
		.din_13 (dout_reg[13]),
		.din_14 (dout_reg[14]),
		.din_15 (dout_reg[15]),
		.din_16 (dout_reg[16]),
		.din_17 (dout_reg[17]),
		.din_18 (dout_reg[18]),
		.din_19 (dout_reg[19]),
		.din_20 (dout_reg[20]),
		.din_21 (dout_reg[21]),
		.din_22 (dout_reg[22]),
		.din_23 (dout_reg[23]),
		.din_24 (dout_reg[24]),
		.din_25 (dout_reg[25]),
		.din_26 (dout_reg[26]),
		.din_27 (dout_reg[27]),
		.din_28 (dout_reg[28]),
		.din_29 (dout_reg[29]),
		.din_30 (dout_reg[30]),
		.din_31 (dout_reg[31]),
		.din_32 (dout_reg[32]),
		.din_33 (dout_reg[33]),
		.din_34 (dout_reg[34]),
		.din_35 (dout_reg[35]),
		.din_36 (dout_reg[36]),
		.din_37 (dout_reg[37]),
		.din_38 (dout_reg[38]),
		.din_39 (dout_reg[39]),
		.din_40 (dout_reg[40]),
		.din_41 (dout_reg[41]),
		.din_42 (dout_reg[42]),
		.din_43 (dout_reg[43]),
		.din_44 (dout_reg[44]),
		.din_45 (dout_reg[45]),
		.din_46 (dout_reg[46]),
		.din_47 (dout_reg[47]),
		.din_48 (dout_reg[48]),
		.din_49 (dout_reg[49]),
		.din_50 (dout_reg[50]),
		.din_51 (dout_reg[51]),
		.din_52 (dout_reg[52]),
		.din_53 (dout_reg[53]),
		.din_54 (dout_reg[54]),
		.din_55 (dout_reg[55]),
		.din_56 (dout_reg[56]),
		.din_57 (dout_reg[57]),
		.din_58 (dout_reg[58]),
		.din_59 (dout_reg[59]),
		.din_60 (dout_reg[60]),
		.din_61 (dout_reg[61]),
		.din_62 (dout_reg[62]),
		.din_63 (dout_reg[63]),
		.din_64 (dout_reg[64]),
		.din_65 (dout_reg[65]),
		.din_66 (dout_reg[66]),
		.din_67 (dout_reg[67]),
		.din_68 (dout_reg[68]),
		.din_69 (dout_reg[69]),
		.din_70 (dout_reg[70]),
		.din_71 (dout_reg[71]),
		.din_72 (dout_reg[72]),
		.din_73 (dout_reg[73]),
		.din_74 (dout_reg[74]),
		.din_75 (dout_reg[75]),
		.din_76 (dout_reg[76]),
		.din_77 (dout_reg[77]),
		.din_78 (dout_reg[78]),
		.din_79 (dout_reg[79]),
		.din_80 (dout_reg[80]),
		.din_81 (dout_reg[81]),
		.din_82 (dout_reg[82]),
		.din_83 (dout_reg[83]),
		.din_84 (dout_reg[84])
	);
endmodule

module reductin_or (
	output wire dout,
	input wire [3:0] din_0,
	input wire [3:0] din_1,
	input wire [3:0] din_2,
	input wire [3:0] din_3,
	input wire [3:0] din_4,
	input wire [3:0] din_5,
	input wire [3:0] din_6,
	input wire [3:0] din_7,
	input wire [3:0] din_8,
	input wire [3:0] din_9,
	input wire [3:0] din_10,
	input wire [3:0] din_11,
	input wire [3:0] din_12,
	input wire [3:0] din_13,
	input wire [3:0] din_14,
	input wire [3:0] din_15,
	input wire [3:0] din_16,
	input wire [3:0] din_17,
	input wire [3:0] din_18,
	input wire [3:0] din_19,
	input wire [3:0] din_20,
	input wire [3:0] din_21,
	input wire [3:0] din_22,
	input wire [3:0] din_23,
	input wire [3:0] din_24,
	input wire [3:0] din_25,
	input wire [3:0] din_26,
	input wire [3:0] din_27,
	input wire [3:0] din_28,
	input wire [3:0] din_29,
	input wire [3:0] din_30,
	input wire [3:0] din_31,
	input wire [3:0] din_32,
	input wire [3:0] din_33,
	input wire [3:0] din_34,
	input wire [3:0] din_35,
	input wire [3:0] din_36,
	input wire [3:0] din_37,
	input wire [3:0] din_38,
	input wire [3:0] din_39,
	input wire [3:0] din_40,
	input wire [3:0] din_41,
	input wire [3:0] din_42,
	input wire [3:0] din_43,
	input wire [3:0] din_44,
	input wire [3:0] din_45,
	input wire [3:0] din_46,
	input wire [3:0] din_47,
	input wire [3:0] din_48,
	input wire [3:0] din_49,
	input wire [3:0] din_50,
	input wire [3:0] din_51,
	input wire [3:0] din_52,
	input wire [3:0] din_53,
	input wire [3:0] din_54,
	input wire [3:0] din_55,
	input wire [3:0] din_56,
	input wire [3:0] din_57,
	input wire [3:0] din_58,
	input wire [3:0] din_59,
	input wire [3:0] din_60,
	input wire [3:0] din_61,
	input wire [3:0] din_62,
	input wire [3:0] din_63,
	input wire [3:0] din_64,
	input wire [3:0] din_65,
	input wire [3:0] din_66,
	input wire [3:0] din_67,
	input wire [3:0] din_68,
	input wire [3:0] din_69,
	input wire [3:0] din_70,
	input wire [3:0] din_71,
	input wire [3:0] din_72,
	input wire [3:0] din_73,
	input wire [3:0] din_74,
	input wire [3:0] din_75,
	input wire [3:0] din_76,
	input wire [3:0] din_77,
	input wire [3:0] din_78,
	input wire [3:0] din_79,
	input wire [3:0] din_80,
	input wire [3:0] din_81,
	input wire [3:0] din_82,
	input wire [3:0] din_83,
	input wire [3:0] din_84
);

assign dout = |{din_0,din_1,din_2,din_3,din_4,din_5,din_6,din_7,din_8,din_9,din_10,din_11,din_12,din_13,din_14,din_15,din_16,din_17,din_18,din_19,din_20,din_21,din_22,din_23,din_24,din_25,din_26,din_27,din_28,din_29,din_30,din_31,din_32,din_33,din_34,din_35,din_36,din_37,din_38,din_39,din_40,din_41,din_42,din_43,din_44,din_45,din_46,din_47,din_48,din_49,din_50,din_51,din_52,din_53,din_54,din_55,din_56,din_57,din_58,din_59,din_60,din_61,din_62,din_63,din_64,din_65,din_66,din_67,din_68,din_69,din_70,din_71,din_72,din_73,din_74,din_75,din_76,din_77,din_78,din_79,din_80,din_81,din_82,din_83,din_84};
endmodule