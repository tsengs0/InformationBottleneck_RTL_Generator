module qsn_left (
	output wire [253:0] sw_out,

	input wire [254:0] sw_in,
	input wire [7:0] sel,
	input wire sys_clk,
	input wire rstn
);

	// Multiplexer Stage 7
	wire [126:0] mux_stage_7;
	assign mux_stage_7[0] = (sel[7] == 1'b1) ? sw_in[128] : sw_in[0];
	assign mux_stage_7[1] = (sel[7] == 1'b1) ? sw_in[129] : sw_in[1];
	assign mux_stage_7[2] = (sel[7] == 1'b1) ? sw_in[130] : sw_in[2];
	assign mux_stage_7[3] = (sel[7] == 1'b1) ? sw_in[131] : sw_in[3];
	assign mux_stage_7[4] = (sel[7] == 1'b1) ? sw_in[132] : sw_in[4];
	assign mux_stage_7[5] = (sel[7] == 1'b1) ? sw_in[133] : sw_in[5];
	assign mux_stage_7[6] = (sel[7] == 1'b1) ? sw_in[134] : sw_in[6];
	assign mux_stage_7[7] = (sel[7] == 1'b1) ? sw_in[135] : sw_in[7];
	assign mux_stage_7[8] = (sel[7] == 1'b1) ? sw_in[136] : sw_in[8];
	assign mux_stage_7[9] = (sel[7] == 1'b1) ? sw_in[137] : sw_in[9];
	assign mux_stage_7[10] = (sel[7] == 1'b1) ? sw_in[138] : sw_in[10];
	assign mux_stage_7[11] = (sel[7] == 1'b1) ? sw_in[139] : sw_in[11];
	assign mux_stage_7[12] = (sel[7] == 1'b1) ? sw_in[140] : sw_in[12];
	assign mux_stage_7[13] = (sel[7] == 1'b1) ? sw_in[141] : sw_in[13];
	assign mux_stage_7[14] = (sel[7] == 1'b1) ? sw_in[142] : sw_in[14];
	assign mux_stage_7[15] = (sel[7] == 1'b1) ? sw_in[143] : sw_in[15];
	assign mux_stage_7[16] = (sel[7] == 1'b1) ? sw_in[144] : sw_in[16];
	assign mux_stage_7[17] = (sel[7] == 1'b1) ? sw_in[145] : sw_in[17];
	assign mux_stage_7[18] = (sel[7] == 1'b1) ? sw_in[146] : sw_in[18];
	assign mux_stage_7[19] = (sel[7] == 1'b1) ? sw_in[147] : sw_in[19];
	assign mux_stage_7[20] = (sel[7] == 1'b1) ? sw_in[148] : sw_in[20];
	assign mux_stage_7[21] = (sel[7] == 1'b1) ? sw_in[149] : sw_in[21];
	assign mux_stage_7[22] = (sel[7] == 1'b1) ? sw_in[150] : sw_in[22];
	assign mux_stage_7[23] = (sel[7] == 1'b1) ? sw_in[151] : sw_in[23];
	assign mux_stage_7[24] = (sel[7] == 1'b1) ? sw_in[152] : sw_in[24];
	assign mux_stage_7[25] = (sel[7] == 1'b1) ? sw_in[153] : sw_in[25];
	assign mux_stage_7[26] = (sel[7] == 1'b1) ? sw_in[154] : sw_in[26];
	assign mux_stage_7[27] = (sel[7] == 1'b1) ? sw_in[155] : sw_in[27];
	assign mux_stage_7[28] = (sel[7] == 1'b1) ? sw_in[156] : sw_in[28];
	assign mux_stage_7[29] = (sel[7] == 1'b1) ? sw_in[157] : sw_in[29];
	assign mux_stage_7[30] = (sel[7] == 1'b1) ? sw_in[158] : sw_in[30];
	assign mux_stage_7[31] = (sel[7] == 1'b1) ? sw_in[159] : sw_in[31];
	assign mux_stage_7[32] = (sel[7] == 1'b1) ? sw_in[160] : sw_in[32];
	assign mux_stage_7[33] = (sel[7] == 1'b1) ? sw_in[161] : sw_in[33];
	assign mux_stage_7[34] = (sel[7] == 1'b1) ? sw_in[162] : sw_in[34];
	assign mux_stage_7[35] = (sel[7] == 1'b1) ? sw_in[163] : sw_in[35];
	assign mux_stage_7[36] = (sel[7] == 1'b1) ? sw_in[164] : sw_in[36];
	assign mux_stage_7[37] = (sel[7] == 1'b1) ? sw_in[165] : sw_in[37];
	assign mux_stage_7[38] = (sel[7] == 1'b1) ? sw_in[166] : sw_in[38];
	assign mux_stage_7[39] = (sel[7] == 1'b1) ? sw_in[167] : sw_in[39];
	assign mux_stage_7[40] = (sel[7] == 1'b1) ? sw_in[168] : sw_in[40];
	assign mux_stage_7[41] = (sel[7] == 1'b1) ? sw_in[169] : sw_in[41];
	assign mux_stage_7[42] = (sel[7] == 1'b1) ? sw_in[170] : sw_in[42];
	assign mux_stage_7[43] = (sel[7] == 1'b1) ? sw_in[171] : sw_in[43];
	assign mux_stage_7[44] = (sel[7] == 1'b1) ? sw_in[172] : sw_in[44];
	assign mux_stage_7[45] = (sel[7] == 1'b1) ? sw_in[173] : sw_in[45];
	assign mux_stage_7[46] = (sel[7] == 1'b1) ? sw_in[174] : sw_in[46];
	assign mux_stage_7[47] = (sel[7] == 1'b1) ? sw_in[175] : sw_in[47];
	assign mux_stage_7[48] = (sel[7] == 1'b1) ? sw_in[176] : sw_in[48];
	assign mux_stage_7[49] = (sel[7] == 1'b1) ? sw_in[177] : sw_in[49];
	assign mux_stage_7[50] = (sel[7] == 1'b1) ? sw_in[178] : sw_in[50];
	assign mux_stage_7[51] = (sel[7] == 1'b1) ? sw_in[179] : sw_in[51];
	assign mux_stage_7[52] = (sel[7] == 1'b1) ? sw_in[180] : sw_in[52];
	assign mux_stage_7[53] = (sel[7] == 1'b1) ? sw_in[181] : sw_in[53];
	assign mux_stage_7[54] = (sel[7] == 1'b1) ? sw_in[182] : sw_in[54];
	assign mux_stage_7[55] = (sel[7] == 1'b1) ? sw_in[183] : sw_in[55];
	assign mux_stage_7[56] = (sel[7] == 1'b1) ? sw_in[184] : sw_in[56];
	assign mux_stage_7[57] = (sel[7] == 1'b1) ? sw_in[185] : sw_in[57];
	assign mux_stage_7[58] = (sel[7] == 1'b1) ? sw_in[186] : sw_in[58];
	assign mux_stage_7[59] = (sel[7] == 1'b1) ? sw_in[187] : sw_in[59];
	assign mux_stage_7[60] = (sel[7] == 1'b1) ? sw_in[188] : sw_in[60];
	assign mux_stage_7[61] = (sel[7] == 1'b1) ? sw_in[189] : sw_in[61];
	assign mux_stage_7[62] = (sel[7] == 1'b1) ? sw_in[190] : sw_in[62];
	assign mux_stage_7[63] = (sel[7] == 1'b1) ? sw_in[191] : sw_in[63];
	assign mux_stage_7[64] = (sel[7] == 1'b1) ? sw_in[192] : sw_in[64];
	assign mux_stage_7[65] = (sel[7] == 1'b1) ? sw_in[193] : sw_in[65];
	assign mux_stage_7[66] = (sel[7] == 1'b1) ? sw_in[194] : sw_in[66];
	assign mux_stage_7[67] = (sel[7] == 1'b1) ? sw_in[195] : sw_in[67];
	assign mux_stage_7[68] = (sel[7] == 1'b1) ? sw_in[196] : sw_in[68];
	assign mux_stage_7[69] = (sel[7] == 1'b1) ? sw_in[197] : sw_in[69];
	assign mux_stage_7[70] = (sel[7] == 1'b1) ? sw_in[198] : sw_in[70];
	assign mux_stage_7[71] = (sel[7] == 1'b1) ? sw_in[199] : sw_in[71];
	assign mux_stage_7[72] = (sel[7] == 1'b1) ? sw_in[200] : sw_in[72];
	assign mux_stage_7[73] = (sel[7] == 1'b1) ? sw_in[201] : sw_in[73];
	assign mux_stage_7[74] = (sel[7] == 1'b1) ? sw_in[202] : sw_in[74];
	assign mux_stage_7[75] = (sel[7] == 1'b1) ? sw_in[203] : sw_in[75];
	assign mux_stage_7[76] = (sel[7] == 1'b1) ? sw_in[204] : sw_in[76];
	assign mux_stage_7[77] = (sel[7] == 1'b1) ? sw_in[205] : sw_in[77];
	assign mux_stage_7[78] = (sel[7] == 1'b1) ? sw_in[206] : sw_in[78];
	assign mux_stage_7[79] = (sel[7] == 1'b1) ? sw_in[207] : sw_in[79];
	assign mux_stage_7[80] = (sel[7] == 1'b1) ? sw_in[208] : sw_in[80];
	assign mux_stage_7[81] = (sel[7] == 1'b1) ? sw_in[209] : sw_in[81];
	assign mux_stage_7[82] = (sel[7] == 1'b1) ? sw_in[210] : sw_in[82];
	assign mux_stage_7[83] = (sel[7] == 1'b1) ? sw_in[211] : sw_in[83];
	assign mux_stage_7[84] = (sel[7] == 1'b1) ? sw_in[212] : sw_in[84];
	assign mux_stage_7[85] = (sel[7] == 1'b1) ? sw_in[213] : sw_in[85];
	assign mux_stage_7[86] = (sel[7] == 1'b1) ? sw_in[214] : sw_in[86];
	assign mux_stage_7[87] = (sel[7] == 1'b1) ? sw_in[215] : sw_in[87];
	assign mux_stage_7[88] = (sel[7] == 1'b1) ? sw_in[216] : sw_in[88];
	assign mux_stage_7[89] = (sel[7] == 1'b1) ? sw_in[217] : sw_in[89];
	assign mux_stage_7[90] = (sel[7] == 1'b1) ? sw_in[218] : sw_in[90];
	assign mux_stage_7[91] = (sel[7] == 1'b1) ? sw_in[219] : sw_in[91];
	assign mux_stage_7[92] = (sel[7] == 1'b1) ? sw_in[220] : sw_in[92];
	assign mux_stage_7[93] = (sel[7] == 1'b1) ? sw_in[221] : sw_in[93];
	assign mux_stage_7[94] = (sel[7] == 1'b1) ? sw_in[222] : sw_in[94];
	assign mux_stage_7[95] = (sel[7] == 1'b1) ? sw_in[223] : sw_in[95];
	assign mux_stage_7[96] = (sel[7] == 1'b1) ? sw_in[224] : sw_in[96];
	assign mux_stage_7[97] = (sel[7] == 1'b1) ? sw_in[225] : sw_in[97];
	assign mux_stage_7[98] = (sel[7] == 1'b1) ? sw_in[226] : sw_in[98];
	assign mux_stage_7[99] = (sel[7] == 1'b1) ? sw_in[227] : sw_in[99];
	assign mux_stage_7[100] = (sel[7] == 1'b1) ? sw_in[228] : sw_in[100];
	assign mux_stage_7[101] = (sel[7] == 1'b1) ? sw_in[229] : sw_in[101];
	assign mux_stage_7[102] = (sel[7] == 1'b1) ? sw_in[230] : sw_in[102];
	assign mux_stage_7[103] = (sel[7] == 1'b1) ? sw_in[231] : sw_in[103];
	assign mux_stage_7[104] = (sel[7] == 1'b1) ? sw_in[232] : sw_in[104];
	assign mux_stage_7[105] = (sel[7] == 1'b1) ? sw_in[233] : sw_in[105];
	assign mux_stage_7[106] = (sel[7] == 1'b1) ? sw_in[234] : sw_in[106];
	assign mux_stage_7[107] = (sel[7] == 1'b1) ? sw_in[235] : sw_in[107];
	assign mux_stage_7[108] = (sel[7] == 1'b1) ? sw_in[236] : sw_in[108];
	assign mux_stage_7[109] = (sel[7] == 1'b1) ? sw_in[237] : sw_in[109];
	assign mux_stage_7[110] = (sel[7] == 1'b1) ? sw_in[238] : sw_in[110];
	assign mux_stage_7[111] = (sel[7] == 1'b1) ? sw_in[239] : sw_in[111];
	assign mux_stage_7[112] = (sel[7] == 1'b1) ? sw_in[240] : sw_in[112];
	assign mux_stage_7[113] = (sel[7] == 1'b1) ? sw_in[241] : sw_in[113];
	assign mux_stage_7[114] = (sel[7] == 1'b1) ? sw_in[242] : sw_in[114];
	assign mux_stage_7[115] = (sel[7] == 1'b1) ? sw_in[243] : sw_in[115];
	assign mux_stage_7[116] = (sel[7] == 1'b1) ? sw_in[244] : sw_in[116];
	assign mux_stage_7[117] = (sel[7] == 1'b1) ? sw_in[245] : sw_in[117];
	assign mux_stage_7[118] = (sel[7] == 1'b1) ? sw_in[246] : sw_in[118];
	assign mux_stage_7[119] = (sel[7] == 1'b1) ? sw_in[247] : sw_in[119];
	assign mux_stage_7[120] = (sel[7] == 1'b1) ? sw_in[248] : sw_in[120];
	assign mux_stage_7[121] = (sel[7] == 1'b1) ? sw_in[249] : sw_in[121];
	assign mux_stage_7[122] = (sel[7] == 1'b1) ? sw_in[250] : sw_in[122];
	assign mux_stage_7[123] = (sel[7] == 1'b1) ? sw_in[251] : sw_in[123];
	assign mux_stage_7[124] = (sel[7] == 1'b1) ? sw_in[252] : sw_in[124];
	assign mux_stage_7[125] = (sel[7] == 1'b1) ? sw_in[253] : sw_in[125];
	assign mux_stage_7[126] = (sel[7] == 1'b1) ? sw_in[254] : sw_in[126];

	// Multiplexer Stage 6
	wire [190:0] mux_stage_6;
	assign mux_stage_6[0] = (sel[6] == 1'b1) ? mux_stage_7[64] : mux_stage_7[0];
	assign mux_stage_6[1] = (sel[6] == 1'b1) ? mux_stage_7[65] : mux_stage_7[1];
	assign mux_stage_6[2] = (sel[6] == 1'b1) ? mux_stage_7[66] : mux_stage_7[2];
	assign mux_stage_6[3] = (sel[6] == 1'b1) ? mux_stage_7[67] : mux_stage_7[3];
	assign mux_stage_6[4] = (sel[6] == 1'b1) ? mux_stage_7[68] : mux_stage_7[4];
	assign mux_stage_6[5] = (sel[6] == 1'b1) ? mux_stage_7[69] : mux_stage_7[5];
	assign mux_stage_6[6] = (sel[6] == 1'b1) ? mux_stage_7[70] : mux_stage_7[6];
	assign mux_stage_6[7] = (sel[6] == 1'b1) ? mux_stage_7[71] : mux_stage_7[7];
	assign mux_stage_6[8] = (sel[6] == 1'b1) ? mux_stage_7[72] : mux_stage_7[8];
	assign mux_stage_6[9] = (sel[6] == 1'b1) ? mux_stage_7[73] : mux_stage_7[9];
	assign mux_stage_6[10] = (sel[6] == 1'b1) ? mux_stage_7[74] : mux_stage_7[10];
	assign mux_stage_6[11] = (sel[6] == 1'b1) ? mux_stage_7[75] : mux_stage_7[11];
	assign mux_stage_6[12] = (sel[6] == 1'b1) ? mux_stage_7[76] : mux_stage_7[12];
	assign mux_stage_6[13] = (sel[6] == 1'b1) ? mux_stage_7[77] : mux_stage_7[13];
	assign mux_stage_6[14] = (sel[6] == 1'b1) ? mux_stage_7[78] : mux_stage_7[14];
	assign mux_stage_6[15] = (sel[6] == 1'b1) ? mux_stage_7[79] : mux_stage_7[15];
	assign mux_stage_6[16] = (sel[6] == 1'b1) ? mux_stage_7[80] : mux_stage_7[16];
	assign mux_stage_6[17] = (sel[6] == 1'b1) ? mux_stage_7[81] : mux_stage_7[17];
	assign mux_stage_6[18] = (sel[6] == 1'b1) ? mux_stage_7[82] : mux_stage_7[18];
	assign mux_stage_6[19] = (sel[6] == 1'b1) ? mux_stage_7[83] : mux_stage_7[19];
	assign mux_stage_6[20] = (sel[6] == 1'b1) ? mux_stage_7[84] : mux_stage_7[20];
	assign mux_stage_6[21] = (sel[6] == 1'b1) ? mux_stage_7[85] : mux_stage_7[21];
	assign mux_stage_6[22] = (sel[6] == 1'b1) ? mux_stage_7[86] : mux_stage_7[22];
	assign mux_stage_6[23] = (sel[6] == 1'b1) ? mux_stage_7[87] : mux_stage_7[23];
	assign mux_stage_6[24] = (sel[6] == 1'b1) ? mux_stage_7[88] : mux_stage_7[24];
	assign mux_stage_6[25] = (sel[6] == 1'b1) ? mux_stage_7[89] : mux_stage_7[25];
	assign mux_stage_6[26] = (sel[6] == 1'b1) ? mux_stage_7[90] : mux_stage_7[26];
	assign mux_stage_6[27] = (sel[6] == 1'b1) ? mux_stage_7[91] : mux_stage_7[27];
	assign mux_stage_6[28] = (sel[6] == 1'b1) ? mux_stage_7[92] : mux_stage_7[28];
	assign mux_stage_6[29] = (sel[6] == 1'b1) ? mux_stage_7[93] : mux_stage_7[29];
	assign mux_stage_6[30] = (sel[6] == 1'b1) ? mux_stage_7[94] : mux_stage_7[30];
	assign mux_stage_6[31] = (sel[6] == 1'b1) ? mux_stage_7[95] : mux_stage_7[31];
	assign mux_stage_6[32] = (sel[6] == 1'b1) ? mux_stage_7[96] : mux_stage_7[32];
	assign mux_stage_6[33] = (sel[6] == 1'b1) ? mux_stage_7[97] : mux_stage_7[33];
	assign mux_stage_6[34] = (sel[6] == 1'b1) ? mux_stage_7[98] : mux_stage_7[34];
	assign mux_stage_6[35] = (sel[6] == 1'b1) ? mux_stage_7[99] : mux_stage_7[35];
	assign mux_stage_6[36] = (sel[6] == 1'b1) ? mux_stage_7[100] : mux_stage_7[36];
	assign mux_stage_6[37] = (sel[6] == 1'b1) ? mux_stage_7[101] : mux_stage_7[37];
	assign mux_stage_6[38] = (sel[6] == 1'b1) ? mux_stage_7[102] : mux_stage_7[38];
	assign mux_stage_6[39] = (sel[6] == 1'b1) ? mux_stage_7[103] : mux_stage_7[39];
	assign mux_stage_6[40] = (sel[6] == 1'b1) ? mux_stage_7[104] : mux_stage_7[40];
	assign mux_stage_6[41] = (sel[6] == 1'b1) ? mux_stage_7[105] : mux_stage_7[41];
	assign mux_stage_6[42] = (sel[6] == 1'b1) ? mux_stage_7[106] : mux_stage_7[42];
	assign mux_stage_6[43] = (sel[6] == 1'b1) ? mux_stage_7[107] : mux_stage_7[43];
	assign mux_stage_6[44] = (sel[6] == 1'b1) ? mux_stage_7[108] : mux_stage_7[44];
	assign mux_stage_6[45] = (sel[6] == 1'b1) ? mux_stage_7[109] : mux_stage_7[45];
	assign mux_stage_6[46] = (sel[6] == 1'b1) ? mux_stage_7[110] : mux_stage_7[46];
	assign mux_stage_6[47] = (sel[6] == 1'b1) ? mux_stage_7[111] : mux_stage_7[47];
	assign mux_stage_6[48] = (sel[6] == 1'b1) ? mux_stage_7[112] : mux_stage_7[48];
	assign mux_stage_6[49] = (sel[6] == 1'b1) ? mux_stage_7[113] : mux_stage_7[49];
	assign mux_stage_6[50] = (sel[6] == 1'b1) ? mux_stage_7[114] : mux_stage_7[50];
	assign mux_stage_6[51] = (sel[6] == 1'b1) ? mux_stage_7[115] : mux_stage_7[51];
	assign mux_stage_6[52] = (sel[6] == 1'b1) ? mux_stage_7[116] : mux_stage_7[52];
	assign mux_stage_6[53] = (sel[6] == 1'b1) ? mux_stage_7[117] : mux_stage_7[53];
	assign mux_stage_6[54] = (sel[6] == 1'b1) ? mux_stage_7[118] : mux_stage_7[54];
	assign mux_stage_6[55] = (sel[6] == 1'b1) ? mux_stage_7[119] : mux_stage_7[55];
	assign mux_stage_6[56] = (sel[6] == 1'b1) ? mux_stage_7[120] : mux_stage_7[56];
	assign mux_stage_6[57] = (sel[6] == 1'b1) ? mux_stage_7[121] : mux_stage_7[57];
	assign mux_stage_6[58] = (sel[6] == 1'b1) ? mux_stage_7[122] : mux_stage_7[58];
	assign mux_stage_6[59] = (sel[6] == 1'b1) ? mux_stage_7[123] : mux_stage_7[59];
	assign mux_stage_6[60] = (sel[6] == 1'b1) ? mux_stage_7[124] : mux_stage_7[60];
	assign mux_stage_6[61] = (sel[6] == 1'b1) ? mux_stage_7[125] : mux_stage_7[61];
	assign mux_stage_6[62] = (sel[6] == 1'b1) ? mux_stage_7[126] : mux_stage_7[62];
	assign mux_stage_6[63] = (sel[6] == 1'b1) ? sw_in[127] : mux_stage_7[63];
	assign mux_stage_6[64] = (sel[6] == 1'b1) ? sw_in[128] : mux_stage_7[64];
	assign mux_stage_6[65] = (sel[6] == 1'b1) ? sw_in[129] : mux_stage_7[65];
	assign mux_stage_6[66] = (sel[6] == 1'b1) ? sw_in[130] : mux_stage_7[66];
	assign mux_stage_6[67] = (sel[6] == 1'b1) ? sw_in[131] : mux_stage_7[67];
	assign mux_stage_6[68] = (sel[6] == 1'b1) ? sw_in[132] : mux_stage_7[68];
	assign mux_stage_6[69] = (sel[6] == 1'b1) ? sw_in[133] : mux_stage_7[69];
	assign mux_stage_6[70] = (sel[6] == 1'b1) ? sw_in[134] : mux_stage_7[70];
	assign mux_stage_6[71] = (sel[6] == 1'b1) ? sw_in[135] : mux_stage_7[71];
	assign mux_stage_6[72] = (sel[6] == 1'b1) ? sw_in[136] : mux_stage_7[72];
	assign mux_stage_6[73] = (sel[6] == 1'b1) ? sw_in[137] : mux_stage_7[73];
	assign mux_stage_6[74] = (sel[6] == 1'b1) ? sw_in[138] : mux_stage_7[74];
	assign mux_stage_6[75] = (sel[6] == 1'b1) ? sw_in[139] : mux_stage_7[75];
	assign mux_stage_6[76] = (sel[6] == 1'b1) ? sw_in[140] : mux_stage_7[76];
	assign mux_stage_6[77] = (sel[6] == 1'b1) ? sw_in[141] : mux_stage_7[77];
	assign mux_stage_6[78] = (sel[6] == 1'b1) ? sw_in[142] : mux_stage_7[78];
	assign mux_stage_6[79] = (sel[6] == 1'b1) ? sw_in[143] : mux_stage_7[79];
	assign mux_stage_6[80] = (sel[6] == 1'b1) ? sw_in[144] : mux_stage_7[80];
	assign mux_stage_6[81] = (sel[6] == 1'b1) ? sw_in[145] : mux_stage_7[81];
	assign mux_stage_6[82] = (sel[6] == 1'b1) ? sw_in[146] : mux_stage_7[82];
	assign mux_stage_6[83] = (sel[6] == 1'b1) ? sw_in[147] : mux_stage_7[83];
	assign mux_stage_6[84] = (sel[6] == 1'b1) ? sw_in[148] : mux_stage_7[84];
	assign mux_stage_6[85] = (sel[6] == 1'b1) ? sw_in[149] : mux_stage_7[85];
	assign mux_stage_6[86] = (sel[6] == 1'b1) ? sw_in[150] : mux_stage_7[86];
	assign mux_stage_6[87] = (sel[6] == 1'b1) ? sw_in[151] : mux_stage_7[87];
	assign mux_stage_6[88] = (sel[6] == 1'b1) ? sw_in[152] : mux_stage_7[88];
	assign mux_stage_6[89] = (sel[6] == 1'b1) ? sw_in[153] : mux_stage_7[89];
	assign mux_stage_6[90] = (sel[6] == 1'b1) ? sw_in[154] : mux_stage_7[90];
	assign mux_stage_6[91] = (sel[6] == 1'b1) ? sw_in[155] : mux_stage_7[91];
	assign mux_stage_6[92] = (sel[6] == 1'b1) ? sw_in[156] : mux_stage_7[92];
	assign mux_stage_6[93] = (sel[6] == 1'b1) ? sw_in[157] : mux_stage_7[93];
	assign mux_stage_6[94] = (sel[6] == 1'b1) ? sw_in[158] : mux_stage_7[94];
	assign mux_stage_6[95] = (sel[6] == 1'b1) ? sw_in[159] : mux_stage_7[95];
	assign mux_stage_6[96] = (sel[6] == 1'b1) ? sw_in[160] : mux_stage_7[96];
	assign mux_stage_6[97] = (sel[6] == 1'b1) ? sw_in[161] : mux_stage_7[97];
	assign mux_stage_6[98] = (sel[6] == 1'b1) ? sw_in[162] : mux_stage_7[98];
	assign mux_stage_6[99] = (sel[6] == 1'b1) ? sw_in[163] : mux_stage_7[99];
	assign mux_stage_6[100] = (sel[6] == 1'b1) ? sw_in[164] : mux_stage_7[100];
	assign mux_stage_6[101] = (sel[6] == 1'b1) ? sw_in[165] : mux_stage_7[101];
	assign mux_stage_6[102] = (sel[6] == 1'b1) ? sw_in[166] : mux_stage_7[102];
	assign mux_stage_6[103] = (sel[6] == 1'b1) ? sw_in[167] : mux_stage_7[103];
	assign mux_stage_6[104] = (sel[6] == 1'b1) ? sw_in[168] : mux_stage_7[104];
	assign mux_stage_6[105] = (sel[6] == 1'b1) ? sw_in[169] : mux_stage_7[105];
	assign mux_stage_6[106] = (sel[6] == 1'b1) ? sw_in[170] : mux_stage_7[106];
	assign mux_stage_6[107] = (sel[6] == 1'b1) ? sw_in[171] : mux_stage_7[107];
	assign mux_stage_6[108] = (sel[6] == 1'b1) ? sw_in[172] : mux_stage_7[108];
	assign mux_stage_6[109] = (sel[6] == 1'b1) ? sw_in[173] : mux_stage_7[109];
	assign mux_stage_6[110] = (sel[6] == 1'b1) ? sw_in[174] : mux_stage_7[110];
	assign mux_stage_6[111] = (sel[6] == 1'b1) ? sw_in[175] : mux_stage_7[111];
	assign mux_stage_6[112] = (sel[6] == 1'b1) ? sw_in[176] : mux_stage_7[112];
	assign mux_stage_6[113] = (sel[6] == 1'b1) ? sw_in[177] : mux_stage_7[113];
	assign mux_stage_6[114] = (sel[6] == 1'b1) ? sw_in[178] : mux_stage_7[114];
	assign mux_stage_6[115] = (sel[6] == 1'b1) ? sw_in[179] : mux_stage_7[115];
	assign mux_stage_6[116] = (sel[6] == 1'b1) ? sw_in[180] : mux_stage_7[116];
	assign mux_stage_6[117] = (sel[6] == 1'b1) ? sw_in[181] : mux_stage_7[117];
	assign mux_stage_6[118] = (sel[6] == 1'b1) ? sw_in[182] : mux_stage_7[118];
	assign mux_stage_6[119] = (sel[6] == 1'b1) ? sw_in[183] : mux_stage_7[119];
	assign mux_stage_6[120] = (sel[6] == 1'b1) ? sw_in[184] : mux_stage_7[120];
	assign mux_stage_6[121] = (sel[6] == 1'b1) ? sw_in[185] : mux_stage_7[121];
	assign mux_stage_6[122] = (sel[6] == 1'b1) ? sw_in[186] : mux_stage_7[122];
	assign mux_stage_6[123] = (sel[6] == 1'b1) ? sw_in[187] : mux_stage_7[123];
	assign mux_stage_6[124] = (sel[6] == 1'b1) ? sw_in[188] : mux_stage_7[124];
	assign mux_stage_6[125] = (sel[6] == 1'b1) ? sw_in[189] : mux_stage_7[125];
	assign mux_stage_6[126] = (sel[6] == 1'b1) ? sw_in[190] : mux_stage_7[126];
	assign mux_stage_6[127] = (sel[6] == 1'b1) ? sw_in[191] : sw_in[127];
	assign mux_stage_6[128] = (sel[6] == 1'b1) ? sw_in[192] : sw_in[128];
	assign mux_stage_6[129] = (sel[6] == 1'b1) ? sw_in[193] : sw_in[129];
	assign mux_stage_6[130] = (sel[6] == 1'b1) ? sw_in[194] : sw_in[130];
	assign mux_stage_6[131] = (sel[6] == 1'b1) ? sw_in[195] : sw_in[131];
	assign mux_stage_6[132] = (sel[6] == 1'b1) ? sw_in[196] : sw_in[132];
	assign mux_stage_6[133] = (sel[6] == 1'b1) ? sw_in[197] : sw_in[133];
	assign mux_stage_6[134] = (sel[6] == 1'b1) ? sw_in[198] : sw_in[134];
	assign mux_stage_6[135] = (sel[6] == 1'b1) ? sw_in[199] : sw_in[135];
	assign mux_stage_6[136] = (sel[6] == 1'b1) ? sw_in[200] : sw_in[136];
	assign mux_stage_6[137] = (sel[6] == 1'b1) ? sw_in[201] : sw_in[137];
	assign mux_stage_6[138] = (sel[6] == 1'b1) ? sw_in[202] : sw_in[138];
	assign mux_stage_6[139] = (sel[6] == 1'b1) ? sw_in[203] : sw_in[139];
	assign mux_stage_6[140] = (sel[6] == 1'b1) ? sw_in[204] : sw_in[140];
	assign mux_stage_6[141] = (sel[6] == 1'b1) ? sw_in[205] : sw_in[141];
	assign mux_stage_6[142] = (sel[6] == 1'b1) ? sw_in[206] : sw_in[142];
	assign mux_stage_6[143] = (sel[6] == 1'b1) ? sw_in[207] : sw_in[143];
	assign mux_stage_6[144] = (sel[6] == 1'b1) ? sw_in[208] : sw_in[144];
	assign mux_stage_6[145] = (sel[6] == 1'b1) ? sw_in[209] : sw_in[145];
	assign mux_stage_6[146] = (sel[6] == 1'b1) ? sw_in[210] : sw_in[146];
	assign mux_stage_6[147] = (sel[6] == 1'b1) ? sw_in[211] : sw_in[147];
	assign mux_stage_6[148] = (sel[6] == 1'b1) ? sw_in[212] : sw_in[148];
	assign mux_stage_6[149] = (sel[6] == 1'b1) ? sw_in[213] : sw_in[149];
	assign mux_stage_6[150] = (sel[6] == 1'b1) ? sw_in[214] : sw_in[150];
	assign mux_stage_6[151] = (sel[6] == 1'b1) ? sw_in[215] : sw_in[151];
	assign mux_stage_6[152] = (sel[6] == 1'b1) ? sw_in[216] : sw_in[152];
	assign mux_stage_6[153] = (sel[6] == 1'b1) ? sw_in[217] : sw_in[153];
	assign mux_stage_6[154] = (sel[6] == 1'b1) ? sw_in[218] : sw_in[154];
	assign mux_stage_6[155] = (sel[6] == 1'b1) ? sw_in[219] : sw_in[155];
	assign mux_stage_6[156] = (sel[6] == 1'b1) ? sw_in[220] : sw_in[156];
	assign mux_stage_6[157] = (sel[6] == 1'b1) ? sw_in[221] : sw_in[157];
	assign mux_stage_6[158] = (sel[6] == 1'b1) ? sw_in[222] : sw_in[158];
	assign mux_stage_6[159] = (sel[6] == 1'b1) ? sw_in[223] : sw_in[159];
	assign mux_stage_6[160] = (sel[6] == 1'b1) ? sw_in[224] : sw_in[160];
	assign mux_stage_6[161] = (sel[6] == 1'b1) ? sw_in[225] : sw_in[161];
	assign mux_stage_6[162] = (sel[6] == 1'b1) ? sw_in[226] : sw_in[162];
	assign mux_stage_6[163] = (sel[6] == 1'b1) ? sw_in[227] : sw_in[163];
	assign mux_stage_6[164] = (sel[6] == 1'b1) ? sw_in[228] : sw_in[164];
	assign mux_stage_6[165] = (sel[6] == 1'b1) ? sw_in[229] : sw_in[165];
	assign mux_stage_6[166] = (sel[6] == 1'b1) ? sw_in[230] : sw_in[166];
	assign mux_stage_6[167] = (sel[6] == 1'b1) ? sw_in[231] : sw_in[167];
	assign mux_stage_6[168] = (sel[6] == 1'b1) ? sw_in[232] : sw_in[168];
	assign mux_stage_6[169] = (sel[6] == 1'b1) ? sw_in[233] : sw_in[169];
	assign mux_stage_6[170] = (sel[6] == 1'b1) ? sw_in[234] : sw_in[170];
	assign mux_stage_6[171] = (sel[6] == 1'b1) ? sw_in[235] : sw_in[171];
	assign mux_stage_6[172] = (sel[6] == 1'b1) ? sw_in[236] : sw_in[172];
	assign mux_stage_6[173] = (sel[6] == 1'b1) ? sw_in[237] : sw_in[173];
	assign mux_stage_6[174] = (sel[6] == 1'b1) ? sw_in[238] : sw_in[174];
	assign mux_stage_6[175] = (sel[6] == 1'b1) ? sw_in[239] : sw_in[175];
	assign mux_stage_6[176] = (sel[6] == 1'b1) ? sw_in[240] : sw_in[176];
	assign mux_stage_6[177] = (sel[6] == 1'b1) ? sw_in[241] : sw_in[177];
	assign mux_stage_6[178] = (sel[6] == 1'b1) ? sw_in[242] : sw_in[178];
	assign mux_stage_6[179] = (sel[6] == 1'b1) ? sw_in[243] : sw_in[179];
	assign mux_stage_6[180] = (sel[6] == 1'b1) ? sw_in[244] : sw_in[180];
	assign mux_stage_6[181] = (sel[6] == 1'b1) ? sw_in[245] : sw_in[181];
	assign mux_stage_6[182] = (sel[6] == 1'b1) ? sw_in[246] : sw_in[182];
	assign mux_stage_6[183] = (sel[6] == 1'b1) ? sw_in[247] : sw_in[183];
	assign mux_stage_6[184] = (sel[6] == 1'b1) ? sw_in[248] : sw_in[184];
	assign mux_stage_6[185] = (sel[6] == 1'b1) ? sw_in[249] : sw_in[185];
	assign mux_stage_6[186] = (sel[6] == 1'b1) ? sw_in[250] : sw_in[186];
	assign mux_stage_6[187] = (sel[6] == 1'b1) ? sw_in[251] : sw_in[187];
	assign mux_stage_6[188] = (sel[6] == 1'b1) ? sw_in[252] : sw_in[188];
	assign mux_stage_6[189] = (sel[6] == 1'b1) ? sw_in[253] : sw_in[189];
	assign mux_stage_6[190] = (sel[6] == 1'b1) ? sw_in[254] : sw_in[190];

	// Multiplexer Stage 5
	wire [222:0] mux_stage_5;
	assign mux_stage_5[0] = (sel[5] == 1'b1) ? mux_stage_6[32] : mux_stage_6[0];
	assign mux_stage_5[1] = (sel[5] == 1'b1) ? mux_stage_6[33] : mux_stage_6[1];
	assign mux_stage_5[2] = (sel[5] == 1'b1) ? mux_stage_6[34] : mux_stage_6[2];
	assign mux_stage_5[3] = (sel[5] == 1'b1) ? mux_stage_6[35] : mux_stage_6[3];
	assign mux_stage_5[4] = (sel[5] == 1'b1) ? mux_stage_6[36] : mux_stage_6[4];
	assign mux_stage_5[5] = (sel[5] == 1'b1) ? mux_stage_6[37] : mux_stage_6[5];
	assign mux_stage_5[6] = (sel[5] == 1'b1) ? mux_stage_6[38] : mux_stage_6[6];
	assign mux_stage_5[7] = (sel[5] == 1'b1) ? mux_stage_6[39] : mux_stage_6[7];
	assign mux_stage_5[8] = (sel[5] == 1'b1) ? mux_stage_6[40] : mux_stage_6[8];
	assign mux_stage_5[9] = (sel[5] == 1'b1) ? mux_stage_6[41] : mux_stage_6[9];
	assign mux_stage_5[10] = (sel[5] == 1'b1) ? mux_stage_6[42] : mux_stage_6[10];
	assign mux_stage_5[11] = (sel[5] == 1'b1) ? mux_stage_6[43] : mux_stage_6[11];
	assign mux_stage_5[12] = (sel[5] == 1'b1) ? mux_stage_6[44] : mux_stage_6[12];
	assign mux_stage_5[13] = (sel[5] == 1'b1) ? mux_stage_6[45] : mux_stage_6[13];
	assign mux_stage_5[14] = (sel[5] == 1'b1) ? mux_stage_6[46] : mux_stage_6[14];
	assign mux_stage_5[15] = (sel[5] == 1'b1) ? mux_stage_6[47] : mux_stage_6[15];
	assign mux_stage_5[16] = (sel[5] == 1'b1) ? mux_stage_6[48] : mux_stage_6[16];
	assign mux_stage_5[17] = (sel[5] == 1'b1) ? mux_stage_6[49] : mux_stage_6[17];
	assign mux_stage_5[18] = (sel[5] == 1'b1) ? mux_stage_6[50] : mux_stage_6[18];
	assign mux_stage_5[19] = (sel[5] == 1'b1) ? mux_stage_6[51] : mux_stage_6[19];
	assign mux_stage_5[20] = (sel[5] == 1'b1) ? mux_stage_6[52] : mux_stage_6[20];
	assign mux_stage_5[21] = (sel[5] == 1'b1) ? mux_stage_6[53] : mux_stage_6[21];
	assign mux_stage_5[22] = (sel[5] == 1'b1) ? mux_stage_6[54] : mux_stage_6[22];
	assign mux_stage_5[23] = (sel[5] == 1'b1) ? mux_stage_6[55] : mux_stage_6[23];
	assign mux_stage_5[24] = (sel[5] == 1'b1) ? mux_stage_6[56] : mux_stage_6[24];
	assign mux_stage_5[25] = (sel[5] == 1'b1) ? mux_stage_6[57] : mux_stage_6[25];
	assign mux_stage_5[26] = (sel[5] == 1'b1) ? mux_stage_6[58] : mux_stage_6[26];
	assign mux_stage_5[27] = (sel[5] == 1'b1) ? mux_stage_6[59] : mux_stage_6[27];
	assign mux_stage_5[28] = (sel[5] == 1'b1) ? mux_stage_6[60] : mux_stage_6[28];
	assign mux_stage_5[29] = (sel[5] == 1'b1) ? mux_stage_6[61] : mux_stage_6[29];
	assign mux_stage_5[30] = (sel[5] == 1'b1) ? mux_stage_6[62] : mux_stage_6[30];
	assign mux_stage_5[31] = (sel[5] == 1'b1) ? mux_stage_6[63] : mux_stage_6[31];
	assign mux_stage_5[32] = (sel[5] == 1'b1) ? mux_stage_6[64] : mux_stage_6[32];
	assign mux_stage_5[33] = (sel[5] == 1'b1) ? mux_stage_6[65] : mux_stage_6[33];
	assign mux_stage_5[34] = (sel[5] == 1'b1) ? mux_stage_6[66] : mux_stage_6[34];
	assign mux_stage_5[35] = (sel[5] == 1'b1) ? mux_stage_6[67] : mux_stage_6[35];
	assign mux_stage_5[36] = (sel[5] == 1'b1) ? mux_stage_6[68] : mux_stage_6[36];
	assign mux_stage_5[37] = (sel[5] == 1'b1) ? mux_stage_6[69] : mux_stage_6[37];
	assign mux_stage_5[38] = (sel[5] == 1'b1) ? mux_stage_6[70] : mux_stage_6[38];
	assign mux_stage_5[39] = (sel[5] == 1'b1) ? mux_stage_6[71] : mux_stage_6[39];
	assign mux_stage_5[40] = (sel[5] == 1'b1) ? mux_stage_6[72] : mux_stage_6[40];
	assign mux_stage_5[41] = (sel[5] == 1'b1) ? mux_stage_6[73] : mux_stage_6[41];
	assign mux_stage_5[42] = (sel[5] == 1'b1) ? mux_stage_6[74] : mux_stage_6[42];
	assign mux_stage_5[43] = (sel[5] == 1'b1) ? mux_stage_6[75] : mux_stage_6[43];
	assign mux_stage_5[44] = (sel[5] == 1'b1) ? mux_stage_6[76] : mux_stage_6[44];
	assign mux_stage_5[45] = (sel[5] == 1'b1) ? mux_stage_6[77] : mux_stage_6[45];
	assign mux_stage_5[46] = (sel[5] == 1'b1) ? mux_stage_6[78] : mux_stage_6[46];
	assign mux_stage_5[47] = (sel[5] == 1'b1) ? mux_stage_6[79] : mux_stage_6[47];
	assign mux_stage_5[48] = (sel[5] == 1'b1) ? mux_stage_6[80] : mux_stage_6[48];
	assign mux_stage_5[49] = (sel[5] == 1'b1) ? mux_stage_6[81] : mux_stage_6[49];
	assign mux_stage_5[50] = (sel[5] == 1'b1) ? mux_stage_6[82] : mux_stage_6[50];
	assign mux_stage_5[51] = (sel[5] == 1'b1) ? mux_stage_6[83] : mux_stage_6[51];
	assign mux_stage_5[52] = (sel[5] == 1'b1) ? mux_stage_6[84] : mux_stage_6[52];
	assign mux_stage_5[53] = (sel[5] == 1'b1) ? mux_stage_6[85] : mux_stage_6[53];
	assign mux_stage_5[54] = (sel[5] == 1'b1) ? mux_stage_6[86] : mux_stage_6[54];
	assign mux_stage_5[55] = (sel[5] == 1'b1) ? mux_stage_6[87] : mux_stage_6[55];
	assign mux_stage_5[56] = (sel[5] == 1'b1) ? mux_stage_6[88] : mux_stage_6[56];
	assign mux_stage_5[57] = (sel[5] == 1'b1) ? mux_stage_6[89] : mux_stage_6[57];
	assign mux_stage_5[58] = (sel[5] == 1'b1) ? mux_stage_6[90] : mux_stage_6[58];
	assign mux_stage_5[59] = (sel[5] == 1'b1) ? mux_stage_6[91] : mux_stage_6[59];
	assign mux_stage_5[60] = (sel[5] == 1'b1) ? mux_stage_6[92] : mux_stage_6[60];
	assign mux_stage_5[61] = (sel[5] == 1'b1) ? mux_stage_6[93] : mux_stage_6[61];
	assign mux_stage_5[62] = (sel[5] == 1'b1) ? mux_stage_6[94] : mux_stage_6[62];
	assign mux_stage_5[63] = (sel[5] == 1'b1) ? mux_stage_6[95] : mux_stage_6[63];
	assign mux_stage_5[64] = (sel[5] == 1'b1) ? mux_stage_6[96] : mux_stage_6[64];
	assign mux_stage_5[65] = (sel[5] == 1'b1) ? mux_stage_6[97] : mux_stage_6[65];
	assign mux_stage_5[66] = (sel[5] == 1'b1) ? mux_stage_6[98] : mux_stage_6[66];
	assign mux_stage_5[67] = (sel[5] == 1'b1) ? mux_stage_6[99] : mux_stage_6[67];
	assign mux_stage_5[68] = (sel[5] == 1'b1) ? mux_stage_6[100] : mux_stage_6[68];
	assign mux_stage_5[69] = (sel[5] == 1'b1) ? mux_stage_6[101] : mux_stage_6[69];
	assign mux_stage_5[70] = (sel[5] == 1'b1) ? mux_stage_6[102] : mux_stage_6[70];
	assign mux_stage_5[71] = (sel[5] == 1'b1) ? mux_stage_6[103] : mux_stage_6[71];
	assign mux_stage_5[72] = (sel[5] == 1'b1) ? mux_stage_6[104] : mux_stage_6[72];
	assign mux_stage_5[73] = (sel[5] == 1'b1) ? mux_stage_6[105] : mux_stage_6[73];
	assign mux_stage_5[74] = (sel[5] == 1'b1) ? mux_stage_6[106] : mux_stage_6[74];
	assign mux_stage_5[75] = (sel[5] == 1'b1) ? mux_stage_6[107] : mux_stage_6[75];
	assign mux_stage_5[76] = (sel[5] == 1'b1) ? mux_stage_6[108] : mux_stage_6[76];
	assign mux_stage_5[77] = (sel[5] == 1'b1) ? mux_stage_6[109] : mux_stage_6[77];
	assign mux_stage_5[78] = (sel[5] == 1'b1) ? mux_stage_6[110] : mux_stage_6[78];
	assign mux_stage_5[79] = (sel[5] == 1'b1) ? mux_stage_6[111] : mux_stage_6[79];
	assign mux_stage_5[80] = (sel[5] == 1'b1) ? mux_stage_6[112] : mux_stage_6[80];
	assign mux_stage_5[81] = (sel[5] == 1'b1) ? mux_stage_6[113] : mux_stage_6[81];
	assign mux_stage_5[82] = (sel[5] == 1'b1) ? mux_stage_6[114] : mux_stage_6[82];
	assign mux_stage_5[83] = (sel[5] == 1'b1) ? mux_stage_6[115] : mux_stage_6[83];
	assign mux_stage_5[84] = (sel[5] == 1'b1) ? mux_stage_6[116] : mux_stage_6[84];
	assign mux_stage_5[85] = (sel[5] == 1'b1) ? mux_stage_6[117] : mux_stage_6[85];
	assign mux_stage_5[86] = (sel[5] == 1'b1) ? mux_stage_6[118] : mux_stage_6[86];
	assign mux_stage_5[87] = (sel[5] == 1'b1) ? mux_stage_6[119] : mux_stage_6[87];
	assign mux_stage_5[88] = (sel[5] == 1'b1) ? mux_stage_6[120] : mux_stage_6[88];
	assign mux_stage_5[89] = (sel[5] == 1'b1) ? mux_stage_6[121] : mux_stage_6[89];
	assign mux_stage_5[90] = (sel[5] == 1'b1) ? mux_stage_6[122] : mux_stage_6[90];
	assign mux_stage_5[91] = (sel[5] == 1'b1) ? mux_stage_6[123] : mux_stage_6[91];
	assign mux_stage_5[92] = (sel[5] == 1'b1) ? mux_stage_6[124] : mux_stage_6[92];
	assign mux_stage_5[93] = (sel[5] == 1'b1) ? mux_stage_6[125] : mux_stage_6[93];
	assign mux_stage_5[94] = (sel[5] == 1'b1) ? mux_stage_6[126] : mux_stage_6[94];
	assign mux_stage_5[95] = (sel[5] == 1'b1) ? mux_stage_6[127] : mux_stage_6[95];
	assign mux_stage_5[96] = (sel[5] == 1'b1) ? mux_stage_6[128] : mux_stage_6[96];
	assign mux_stage_5[97] = (sel[5] == 1'b1) ? mux_stage_6[129] : mux_stage_6[97];
	assign mux_stage_5[98] = (sel[5] == 1'b1) ? mux_stage_6[130] : mux_stage_6[98];
	assign mux_stage_5[99] = (sel[5] == 1'b1) ? mux_stage_6[131] : mux_stage_6[99];
	assign mux_stage_5[100] = (sel[5] == 1'b1) ? mux_stage_6[132] : mux_stage_6[100];
	assign mux_stage_5[101] = (sel[5] == 1'b1) ? mux_stage_6[133] : mux_stage_6[101];
	assign mux_stage_5[102] = (sel[5] == 1'b1) ? mux_stage_6[134] : mux_stage_6[102];
	assign mux_stage_5[103] = (sel[5] == 1'b1) ? mux_stage_6[135] : mux_stage_6[103];
	assign mux_stage_5[104] = (sel[5] == 1'b1) ? mux_stage_6[136] : mux_stage_6[104];
	assign mux_stage_5[105] = (sel[5] == 1'b1) ? mux_stage_6[137] : mux_stage_6[105];
	assign mux_stage_5[106] = (sel[5] == 1'b1) ? mux_stage_6[138] : mux_stage_6[106];
	assign mux_stage_5[107] = (sel[5] == 1'b1) ? mux_stage_6[139] : mux_stage_6[107];
	assign mux_stage_5[108] = (sel[5] == 1'b1) ? mux_stage_6[140] : mux_stage_6[108];
	assign mux_stage_5[109] = (sel[5] == 1'b1) ? mux_stage_6[141] : mux_stage_6[109];
	assign mux_stage_5[110] = (sel[5] == 1'b1) ? mux_stage_6[142] : mux_stage_6[110];
	assign mux_stage_5[111] = (sel[5] == 1'b1) ? mux_stage_6[143] : mux_stage_6[111];
	assign mux_stage_5[112] = (sel[5] == 1'b1) ? mux_stage_6[144] : mux_stage_6[112];
	assign mux_stage_5[113] = (sel[5] == 1'b1) ? mux_stage_6[145] : mux_stage_6[113];
	assign mux_stage_5[114] = (sel[5] == 1'b1) ? mux_stage_6[146] : mux_stage_6[114];
	assign mux_stage_5[115] = (sel[5] == 1'b1) ? mux_stage_6[147] : mux_stage_6[115];
	assign mux_stage_5[116] = (sel[5] == 1'b1) ? mux_stage_6[148] : mux_stage_6[116];
	assign mux_stage_5[117] = (sel[5] == 1'b1) ? mux_stage_6[149] : mux_stage_6[117];
	assign mux_stage_5[118] = (sel[5] == 1'b1) ? mux_stage_6[150] : mux_stage_6[118];
	assign mux_stage_5[119] = (sel[5] == 1'b1) ? mux_stage_6[151] : mux_stage_6[119];
	assign mux_stage_5[120] = (sel[5] == 1'b1) ? mux_stage_6[152] : mux_stage_6[120];
	assign mux_stage_5[121] = (sel[5] == 1'b1) ? mux_stage_6[153] : mux_stage_6[121];
	assign mux_stage_5[122] = (sel[5] == 1'b1) ? mux_stage_6[154] : mux_stage_6[122];
	assign mux_stage_5[123] = (sel[5] == 1'b1) ? mux_stage_6[155] : mux_stage_6[123];
	assign mux_stage_5[124] = (sel[5] == 1'b1) ? mux_stage_6[156] : mux_stage_6[124];
	assign mux_stage_5[125] = (sel[5] == 1'b1) ? mux_stage_6[157] : mux_stage_6[125];
	assign mux_stage_5[126] = (sel[5] == 1'b1) ? mux_stage_6[158] : mux_stage_6[126];
	assign mux_stage_5[127] = (sel[5] == 1'b1) ? mux_stage_6[159] : mux_stage_6[127];
	assign mux_stage_5[128] = (sel[5] == 1'b1) ? mux_stage_6[160] : mux_stage_6[128];
	assign mux_stage_5[129] = (sel[5] == 1'b1) ? mux_stage_6[161] : mux_stage_6[129];
	assign mux_stage_5[130] = (sel[5] == 1'b1) ? mux_stage_6[162] : mux_stage_6[130];
	assign mux_stage_5[131] = (sel[5] == 1'b1) ? mux_stage_6[163] : mux_stage_6[131];
	assign mux_stage_5[132] = (sel[5] == 1'b1) ? mux_stage_6[164] : mux_stage_6[132];
	assign mux_stage_5[133] = (sel[5] == 1'b1) ? mux_stage_6[165] : mux_stage_6[133];
	assign mux_stage_5[134] = (sel[5] == 1'b1) ? mux_stage_6[166] : mux_stage_6[134];
	assign mux_stage_5[135] = (sel[5] == 1'b1) ? mux_stage_6[167] : mux_stage_6[135];
	assign mux_stage_5[136] = (sel[5] == 1'b1) ? mux_stage_6[168] : mux_stage_6[136];
	assign mux_stage_5[137] = (sel[5] == 1'b1) ? mux_stage_6[169] : mux_stage_6[137];
	assign mux_stage_5[138] = (sel[5] == 1'b1) ? mux_stage_6[170] : mux_stage_6[138];
	assign mux_stage_5[139] = (sel[5] == 1'b1) ? mux_stage_6[171] : mux_stage_6[139];
	assign mux_stage_5[140] = (sel[5] == 1'b1) ? mux_stage_6[172] : mux_stage_6[140];
	assign mux_stage_5[141] = (sel[5] == 1'b1) ? mux_stage_6[173] : mux_stage_6[141];
	assign mux_stage_5[142] = (sel[5] == 1'b1) ? mux_stage_6[174] : mux_stage_6[142];
	assign mux_stage_5[143] = (sel[5] == 1'b1) ? mux_stage_6[175] : mux_stage_6[143];
	assign mux_stage_5[144] = (sel[5] == 1'b1) ? mux_stage_6[176] : mux_stage_6[144];
	assign mux_stage_5[145] = (sel[5] == 1'b1) ? mux_stage_6[177] : mux_stage_6[145];
	assign mux_stage_5[146] = (sel[5] == 1'b1) ? mux_stage_6[178] : mux_stage_6[146];
	assign mux_stage_5[147] = (sel[5] == 1'b1) ? mux_stage_6[179] : mux_stage_6[147];
	assign mux_stage_5[148] = (sel[5] == 1'b1) ? mux_stage_6[180] : mux_stage_6[148];
	assign mux_stage_5[149] = (sel[5] == 1'b1) ? mux_stage_6[181] : mux_stage_6[149];
	assign mux_stage_5[150] = (sel[5] == 1'b1) ? mux_stage_6[182] : mux_stage_6[150];
	assign mux_stage_5[151] = (sel[5] == 1'b1) ? mux_stage_6[183] : mux_stage_6[151];
	assign mux_stage_5[152] = (sel[5] == 1'b1) ? mux_stage_6[184] : mux_stage_6[152];
	assign mux_stage_5[153] = (sel[5] == 1'b1) ? mux_stage_6[185] : mux_stage_6[153];
	assign mux_stage_5[154] = (sel[5] == 1'b1) ? mux_stage_6[186] : mux_stage_6[154];
	assign mux_stage_5[155] = (sel[5] == 1'b1) ? mux_stage_6[187] : mux_stage_6[155];
	assign mux_stage_5[156] = (sel[5] == 1'b1) ? mux_stage_6[188] : mux_stage_6[156];
	assign mux_stage_5[157] = (sel[5] == 1'b1) ? mux_stage_6[189] : mux_stage_6[157];
	assign mux_stage_5[158] = (sel[5] == 1'b1) ? mux_stage_6[190] : mux_stage_6[158];
	assign mux_stage_5[159] = (sel[5] == 1'b1) ? sw_in[191] : mux_stage_6[159];
	assign mux_stage_5[160] = (sel[5] == 1'b1) ? sw_in[192] : mux_stage_6[160];
	assign mux_stage_5[161] = (sel[5] == 1'b1) ? sw_in[193] : mux_stage_6[161];
	assign mux_stage_5[162] = (sel[5] == 1'b1) ? sw_in[194] : mux_stage_6[162];
	assign mux_stage_5[163] = (sel[5] == 1'b1) ? sw_in[195] : mux_stage_6[163];
	assign mux_stage_5[164] = (sel[5] == 1'b1) ? sw_in[196] : mux_stage_6[164];
	assign mux_stage_5[165] = (sel[5] == 1'b1) ? sw_in[197] : mux_stage_6[165];
	assign mux_stage_5[166] = (sel[5] == 1'b1) ? sw_in[198] : mux_stage_6[166];
	assign mux_stage_5[167] = (sel[5] == 1'b1) ? sw_in[199] : mux_stage_6[167];
	assign mux_stage_5[168] = (sel[5] == 1'b1) ? sw_in[200] : mux_stage_6[168];
	assign mux_stage_5[169] = (sel[5] == 1'b1) ? sw_in[201] : mux_stage_6[169];
	assign mux_stage_5[170] = (sel[5] == 1'b1) ? sw_in[202] : mux_stage_6[170];
	assign mux_stage_5[171] = (sel[5] == 1'b1) ? sw_in[203] : mux_stage_6[171];
	assign mux_stage_5[172] = (sel[5] == 1'b1) ? sw_in[204] : mux_stage_6[172];
	assign mux_stage_5[173] = (sel[5] == 1'b1) ? sw_in[205] : mux_stage_6[173];
	assign mux_stage_5[174] = (sel[5] == 1'b1) ? sw_in[206] : mux_stage_6[174];
	assign mux_stage_5[175] = (sel[5] == 1'b1) ? sw_in[207] : mux_stage_6[175];
	assign mux_stage_5[176] = (sel[5] == 1'b1) ? sw_in[208] : mux_stage_6[176];
	assign mux_stage_5[177] = (sel[5] == 1'b1) ? sw_in[209] : mux_stage_6[177];
	assign mux_stage_5[178] = (sel[5] == 1'b1) ? sw_in[210] : mux_stage_6[178];
	assign mux_stage_5[179] = (sel[5] == 1'b1) ? sw_in[211] : mux_stage_6[179];
	assign mux_stage_5[180] = (sel[5] == 1'b1) ? sw_in[212] : mux_stage_6[180];
	assign mux_stage_5[181] = (sel[5] == 1'b1) ? sw_in[213] : mux_stage_6[181];
	assign mux_stage_5[182] = (sel[5] == 1'b1) ? sw_in[214] : mux_stage_6[182];
	assign mux_stage_5[183] = (sel[5] == 1'b1) ? sw_in[215] : mux_stage_6[183];
	assign mux_stage_5[184] = (sel[5] == 1'b1) ? sw_in[216] : mux_stage_6[184];
	assign mux_stage_5[185] = (sel[5] == 1'b1) ? sw_in[217] : mux_stage_6[185];
	assign mux_stage_5[186] = (sel[5] == 1'b1) ? sw_in[218] : mux_stage_6[186];
	assign mux_stage_5[187] = (sel[5] == 1'b1) ? sw_in[219] : mux_stage_6[187];
	assign mux_stage_5[188] = (sel[5] == 1'b1) ? sw_in[220] : mux_stage_6[188];
	assign mux_stage_5[189] = (sel[5] == 1'b1) ? sw_in[221] : mux_stage_6[189];
	assign mux_stage_5[190] = (sel[5] == 1'b1) ? sw_in[222] : mux_stage_6[190];
	assign mux_stage_5[191] = (sel[5] == 1'b1) ? sw_in[223] : sw_in[191];
	assign mux_stage_5[192] = (sel[5] == 1'b1) ? sw_in[224] : sw_in[192];
	assign mux_stage_5[193] = (sel[5] == 1'b1) ? sw_in[225] : sw_in[193];
	assign mux_stage_5[194] = (sel[5] == 1'b1) ? sw_in[226] : sw_in[194];
	assign mux_stage_5[195] = (sel[5] == 1'b1) ? sw_in[227] : sw_in[195];
	assign mux_stage_5[196] = (sel[5] == 1'b1) ? sw_in[228] : sw_in[196];
	assign mux_stage_5[197] = (sel[5] == 1'b1) ? sw_in[229] : sw_in[197];
	assign mux_stage_5[198] = (sel[5] == 1'b1) ? sw_in[230] : sw_in[198];
	assign mux_stage_5[199] = (sel[5] == 1'b1) ? sw_in[231] : sw_in[199];
	assign mux_stage_5[200] = (sel[5] == 1'b1) ? sw_in[232] : sw_in[200];
	assign mux_stage_5[201] = (sel[5] == 1'b1) ? sw_in[233] : sw_in[201];
	assign mux_stage_5[202] = (sel[5] == 1'b1) ? sw_in[234] : sw_in[202];
	assign mux_stage_5[203] = (sel[5] == 1'b1) ? sw_in[235] : sw_in[203];
	assign mux_stage_5[204] = (sel[5] == 1'b1) ? sw_in[236] : sw_in[204];
	assign mux_stage_5[205] = (sel[5] == 1'b1) ? sw_in[237] : sw_in[205];
	assign mux_stage_5[206] = (sel[5] == 1'b1) ? sw_in[238] : sw_in[206];
	assign mux_stage_5[207] = (sel[5] == 1'b1) ? sw_in[239] : sw_in[207];
	assign mux_stage_5[208] = (sel[5] == 1'b1) ? sw_in[240] : sw_in[208];
	assign mux_stage_5[209] = (sel[5] == 1'b1) ? sw_in[241] : sw_in[209];
	assign mux_stage_5[210] = (sel[5] == 1'b1) ? sw_in[242] : sw_in[210];
	assign mux_stage_5[211] = (sel[5] == 1'b1) ? sw_in[243] : sw_in[211];
	assign mux_stage_5[212] = (sel[5] == 1'b1) ? sw_in[244] : sw_in[212];
	assign mux_stage_5[213] = (sel[5] == 1'b1) ? sw_in[245] : sw_in[213];
	assign mux_stage_5[214] = (sel[5] == 1'b1) ? sw_in[246] : sw_in[214];
	assign mux_stage_5[215] = (sel[5] == 1'b1) ? sw_in[247] : sw_in[215];
	assign mux_stage_5[216] = (sel[5] == 1'b1) ? sw_in[248] : sw_in[216];
	assign mux_stage_5[217] = (sel[5] == 1'b1) ? sw_in[249] : sw_in[217];
	assign mux_stage_5[218] = (sel[5] == 1'b1) ? sw_in[250] : sw_in[218];
	assign mux_stage_5[219] = (sel[5] == 1'b1) ? sw_in[251] : sw_in[219];
	assign mux_stage_5[220] = (sel[5] == 1'b1) ? sw_in[252] : sw_in[220];
	assign mux_stage_5[221] = (sel[5] == 1'b1) ? sw_in[253] : sw_in[221];
	assign mux_stage_5[222] = (sel[5] == 1'b1) ? sw_in[254] : sw_in[222];

	// Multiplexer Stage 4
	reg [238:0] mux_stage_4;
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[0] <= 0; else if(sel[4] == 1'b1) mux_stage_4[0] <= mux_stage_5[16]; else mux_stage_4[0] <= mux_stage_5[0]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[1] <= 0; else if(sel[4] == 1'b1) mux_stage_4[1] <= mux_stage_5[17]; else mux_stage_4[1] <= mux_stage_5[1]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[2] <= 0; else if(sel[4] == 1'b1) mux_stage_4[2] <= mux_stage_5[18]; else mux_stage_4[2] <= mux_stage_5[2]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[3] <= 0; else if(sel[4] == 1'b1) mux_stage_4[3] <= mux_stage_5[19]; else mux_stage_4[3] <= mux_stage_5[3]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[4] <= 0; else if(sel[4] == 1'b1) mux_stage_4[4] <= mux_stage_5[20]; else mux_stage_4[4] <= mux_stage_5[4]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[5] <= 0; else if(sel[4] == 1'b1) mux_stage_4[5] <= mux_stage_5[21]; else mux_stage_4[5] <= mux_stage_5[5]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[6] <= 0; else if(sel[4] == 1'b1) mux_stage_4[6] <= mux_stage_5[22]; else mux_stage_4[6] <= mux_stage_5[6]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[7] <= 0; else if(sel[4] == 1'b1) mux_stage_4[7] <= mux_stage_5[23]; else mux_stage_4[7] <= mux_stage_5[7]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[8] <= 0; else if(sel[4] == 1'b1) mux_stage_4[8] <= mux_stage_5[24]; else mux_stage_4[8] <= mux_stage_5[8]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[9] <= 0; else if(sel[4] == 1'b1) mux_stage_4[9] <= mux_stage_5[25]; else mux_stage_4[9] <= mux_stage_5[9]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[10] <= 0; else if(sel[4] == 1'b1) mux_stage_4[10] <= mux_stage_5[26]; else mux_stage_4[10] <= mux_stage_5[10]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[11] <= 0; else if(sel[4] == 1'b1) mux_stage_4[11] <= mux_stage_5[27]; else mux_stage_4[11] <= mux_stage_5[11]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[12] <= 0; else if(sel[4] == 1'b1) mux_stage_4[12] <= mux_stage_5[28]; else mux_stage_4[12] <= mux_stage_5[12]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[13] <= 0; else if(sel[4] == 1'b1) mux_stage_4[13] <= mux_stage_5[29]; else mux_stage_4[13] <= mux_stage_5[13]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[14] <= 0; else if(sel[4] == 1'b1) mux_stage_4[14] <= mux_stage_5[30]; else mux_stage_4[14] <= mux_stage_5[14]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[15] <= 0; else if(sel[4] == 1'b1) mux_stage_4[15] <= mux_stage_5[31]; else mux_stage_4[15] <= mux_stage_5[15]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[16] <= 0; else if(sel[4] == 1'b1) mux_stage_4[16] <= mux_stage_5[32]; else mux_stage_4[16] <= mux_stage_5[16]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[17] <= 0; else if(sel[4] == 1'b1) mux_stage_4[17] <= mux_stage_5[33]; else mux_stage_4[17] <= mux_stage_5[17]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[18] <= 0; else if(sel[4] == 1'b1) mux_stage_4[18] <= mux_stage_5[34]; else mux_stage_4[18] <= mux_stage_5[18]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[19] <= 0; else if(sel[4] == 1'b1) mux_stage_4[19] <= mux_stage_5[35]; else mux_stage_4[19] <= mux_stage_5[19]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[20] <= 0; else if(sel[4] == 1'b1) mux_stage_4[20] <= mux_stage_5[36]; else mux_stage_4[20] <= mux_stage_5[20]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[21] <= 0; else if(sel[4] == 1'b1) mux_stage_4[21] <= mux_stage_5[37]; else mux_stage_4[21] <= mux_stage_5[21]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[22] <= 0; else if(sel[4] == 1'b1) mux_stage_4[22] <= mux_stage_5[38]; else mux_stage_4[22] <= mux_stage_5[22]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[23] <= 0; else if(sel[4] == 1'b1) mux_stage_4[23] <= mux_stage_5[39]; else mux_stage_4[23] <= mux_stage_5[23]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[24] <= 0; else if(sel[4] == 1'b1) mux_stage_4[24] <= mux_stage_5[40]; else mux_stage_4[24] <= mux_stage_5[24]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[25] <= 0; else if(sel[4] == 1'b1) mux_stage_4[25] <= mux_stage_5[41]; else mux_stage_4[25] <= mux_stage_5[25]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[26] <= 0; else if(sel[4] == 1'b1) mux_stage_4[26] <= mux_stage_5[42]; else mux_stage_4[26] <= mux_stage_5[26]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[27] <= 0; else if(sel[4] == 1'b1) mux_stage_4[27] <= mux_stage_5[43]; else mux_stage_4[27] <= mux_stage_5[27]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[28] <= 0; else if(sel[4] == 1'b1) mux_stage_4[28] <= mux_stage_5[44]; else mux_stage_4[28] <= mux_stage_5[28]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[29] <= 0; else if(sel[4] == 1'b1) mux_stage_4[29] <= mux_stage_5[45]; else mux_stage_4[29] <= mux_stage_5[29]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[30] <= 0; else if(sel[4] == 1'b1) mux_stage_4[30] <= mux_stage_5[46]; else mux_stage_4[30] <= mux_stage_5[30]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[31] <= 0; else if(sel[4] == 1'b1) mux_stage_4[31] <= mux_stage_5[47]; else mux_stage_4[31] <= mux_stage_5[31]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[32] <= 0; else if(sel[4] == 1'b1) mux_stage_4[32] <= mux_stage_5[48]; else mux_stage_4[32] <= mux_stage_5[32]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[33] <= 0; else if(sel[4] == 1'b1) mux_stage_4[33] <= mux_stage_5[49]; else mux_stage_4[33] <= mux_stage_5[33]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[34] <= 0; else if(sel[4] == 1'b1) mux_stage_4[34] <= mux_stage_5[50]; else mux_stage_4[34] <= mux_stage_5[34]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[35] <= 0; else if(sel[4] == 1'b1) mux_stage_4[35] <= mux_stage_5[51]; else mux_stage_4[35] <= mux_stage_5[35]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[36] <= 0; else if(sel[4] == 1'b1) mux_stage_4[36] <= mux_stage_5[52]; else mux_stage_4[36] <= mux_stage_5[36]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[37] <= 0; else if(sel[4] == 1'b1) mux_stage_4[37] <= mux_stage_5[53]; else mux_stage_4[37] <= mux_stage_5[37]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[38] <= 0; else if(sel[4] == 1'b1) mux_stage_4[38] <= mux_stage_5[54]; else mux_stage_4[38] <= mux_stage_5[38]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[39] <= 0; else if(sel[4] == 1'b1) mux_stage_4[39] <= mux_stage_5[55]; else mux_stage_4[39] <= mux_stage_5[39]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[40] <= 0; else if(sel[4] == 1'b1) mux_stage_4[40] <= mux_stage_5[56]; else mux_stage_4[40] <= mux_stage_5[40]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[41] <= 0; else if(sel[4] == 1'b1) mux_stage_4[41] <= mux_stage_5[57]; else mux_stage_4[41] <= mux_stage_5[41]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[42] <= 0; else if(sel[4] == 1'b1) mux_stage_4[42] <= mux_stage_5[58]; else mux_stage_4[42] <= mux_stage_5[42]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[43] <= 0; else if(sel[4] == 1'b1) mux_stage_4[43] <= mux_stage_5[59]; else mux_stage_4[43] <= mux_stage_5[43]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[44] <= 0; else if(sel[4] == 1'b1) mux_stage_4[44] <= mux_stage_5[60]; else mux_stage_4[44] <= mux_stage_5[44]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[45] <= 0; else if(sel[4] == 1'b1) mux_stage_4[45] <= mux_stage_5[61]; else mux_stage_4[45] <= mux_stage_5[45]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[46] <= 0; else if(sel[4] == 1'b1) mux_stage_4[46] <= mux_stage_5[62]; else mux_stage_4[46] <= mux_stage_5[46]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[47] <= 0; else if(sel[4] == 1'b1) mux_stage_4[47] <= mux_stage_5[63]; else mux_stage_4[47] <= mux_stage_5[47]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[48] <= 0; else if(sel[4] == 1'b1) mux_stage_4[48] <= mux_stage_5[64]; else mux_stage_4[48] <= mux_stage_5[48]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[49] <= 0; else if(sel[4] == 1'b1) mux_stage_4[49] <= mux_stage_5[65]; else mux_stage_4[49] <= mux_stage_5[49]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[50] <= 0; else if(sel[4] == 1'b1) mux_stage_4[50] <= mux_stage_5[66]; else mux_stage_4[50] <= mux_stage_5[50]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[51] <= 0; else if(sel[4] == 1'b1) mux_stage_4[51] <= mux_stage_5[67]; else mux_stage_4[51] <= mux_stage_5[51]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[52] <= 0; else if(sel[4] == 1'b1) mux_stage_4[52] <= mux_stage_5[68]; else mux_stage_4[52] <= mux_stage_5[52]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[53] <= 0; else if(sel[4] == 1'b1) mux_stage_4[53] <= mux_stage_5[69]; else mux_stage_4[53] <= mux_stage_5[53]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[54] <= 0; else if(sel[4] == 1'b1) mux_stage_4[54] <= mux_stage_5[70]; else mux_stage_4[54] <= mux_stage_5[54]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[55] <= 0; else if(sel[4] == 1'b1) mux_stage_4[55] <= mux_stage_5[71]; else mux_stage_4[55] <= mux_stage_5[55]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[56] <= 0; else if(sel[4] == 1'b1) mux_stage_4[56] <= mux_stage_5[72]; else mux_stage_4[56] <= mux_stage_5[56]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[57] <= 0; else if(sel[4] == 1'b1) mux_stage_4[57] <= mux_stage_5[73]; else mux_stage_4[57] <= mux_stage_5[57]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[58] <= 0; else if(sel[4] == 1'b1) mux_stage_4[58] <= mux_stage_5[74]; else mux_stage_4[58] <= mux_stage_5[58]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[59] <= 0; else if(sel[4] == 1'b1) mux_stage_4[59] <= mux_stage_5[75]; else mux_stage_4[59] <= mux_stage_5[59]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[60] <= 0; else if(sel[4] == 1'b1) mux_stage_4[60] <= mux_stage_5[76]; else mux_stage_4[60] <= mux_stage_5[60]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[61] <= 0; else if(sel[4] == 1'b1) mux_stage_4[61] <= mux_stage_5[77]; else mux_stage_4[61] <= mux_stage_5[61]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[62] <= 0; else if(sel[4] == 1'b1) mux_stage_4[62] <= mux_stage_5[78]; else mux_stage_4[62] <= mux_stage_5[62]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[63] <= 0; else if(sel[4] == 1'b1) mux_stage_4[63] <= mux_stage_5[79]; else mux_stage_4[63] <= mux_stage_5[63]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[64] <= 0; else if(sel[4] == 1'b1) mux_stage_4[64] <= mux_stage_5[80]; else mux_stage_4[64] <= mux_stage_5[64]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[65] <= 0; else if(sel[4] == 1'b1) mux_stage_4[65] <= mux_stage_5[81]; else mux_stage_4[65] <= mux_stage_5[65]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[66] <= 0; else if(sel[4] == 1'b1) mux_stage_4[66] <= mux_stage_5[82]; else mux_stage_4[66] <= mux_stage_5[66]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[67] <= 0; else if(sel[4] == 1'b1) mux_stage_4[67] <= mux_stage_5[83]; else mux_stage_4[67] <= mux_stage_5[67]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[68] <= 0; else if(sel[4] == 1'b1) mux_stage_4[68] <= mux_stage_5[84]; else mux_stage_4[68] <= mux_stage_5[68]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[69] <= 0; else if(sel[4] == 1'b1) mux_stage_4[69] <= mux_stage_5[85]; else mux_stage_4[69] <= mux_stage_5[69]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[70] <= 0; else if(sel[4] == 1'b1) mux_stage_4[70] <= mux_stage_5[86]; else mux_stage_4[70] <= mux_stage_5[70]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[71] <= 0; else if(sel[4] == 1'b1) mux_stage_4[71] <= mux_stage_5[87]; else mux_stage_4[71] <= mux_stage_5[71]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[72] <= 0; else if(sel[4] == 1'b1) mux_stage_4[72] <= mux_stage_5[88]; else mux_stage_4[72] <= mux_stage_5[72]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[73] <= 0; else if(sel[4] == 1'b1) mux_stage_4[73] <= mux_stage_5[89]; else mux_stage_4[73] <= mux_stage_5[73]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[74] <= 0; else if(sel[4] == 1'b1) mux_stage_4[74] <= mux_stage_5[90]; else mux_stage_4[74] <= mux_stage_5[74]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[75] <= 0; else if(sel[4] == 1'b1) mux_stage_4[75] <= mux_stage_5[91]; else mux_stage_4[75] <= mux_stage_5[75]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[76] <= 0; else if(sel[4] == 1'b1) mux_stage_4[76] <= mux_stage_5[92]; else mux_stage_4[76] <= mux_stage_5[76]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[77] <= 0; else if(sel[4] == 1'b1) mux_stage_4[77] <= mux_stage_5[93]; else mux_stage_4[77] <= mux_stage_5[77]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[78] <= 0; else if(sel[4] == 1'b1) mux_stage_4[78] <= mux_stage_5[94]; else mux_stage_4[78] <= mux_stage_5[78]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[79] <= 0; else if(sel[4] == 1'b1) mux_stage_4[79] <= mux_stage_5[95]; else mux_stage_4[79] <= mux_stage_5[79]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[80] <= 0; else if(sel[4] == 1'b1) mux_stage_4[80] <= mux_stage_5[96]; else mux_stage_4[80] <= mux_stage_5[80]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[81] <= 0; else if(sel[4] == 1'b1) mux_stage_4[81] <= mux_stage_5[97]; else mux_stage_4[81] <= mux_stage_5[81]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[82] <= 0; else if(sel[4] == 1'b1) mux_stage_4[82] <= mux_stage_5[98]; else mux_stage_4[82] <= mux_stage_5[82]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[83] <= 0; else if(sel[4] == 1'b1) mux_stage_4[83] <= mux_stage_5[99]; else mux_stage_4[83] <= mux_stage_5[83]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[84] <= 0; else if(sel[4] == 1'b1) mux_stage_4[84] <= mux_stage_5[100]; else mux_stage_4[84] <= mux_stage_5[84]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[85] <= 0; else if(sel[4] == 1'b1) mux_stage_4[85] <= mux_stage_5[101]; else mux_stage_4[85] <= mux_stage_5[85]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[86] <= 0; else if(sel[4] == 1'b1) mux_stage_4[86] <= mux_stage_5[102]; else mux_stage_4[86] <= mux_stage_5[86]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[87] <= 0; else if(sel[4] == 1'b1) mux_stage_4[87] <= mux_stage_5[103]; else mux_stage_4[87] <= mux_stage_5[87]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[88] <= 0; else if(sel[4] == 1'b1) mux_stage_4[88] <= mux_stage_5[104]; else mux_stage_4[88] <= mux_stage_5[88]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[89] <= 0; else if(sel[4] == 1'b1) mux_stage_4[89] <= mux_stage_5[105]; else mux_stage_4[89] <= mux_stage_5[89]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[90] <= 0; else if(sel[4] == 1'b1) mux_stage_4[90] <= mux_stage_5[106]; else mux_stage_4[90] <= mux_stage_5[90]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[91] <= 0; else if(sel[4] == 1'b1) mux_stage_4[91] <= mux_stage_5[107]; else mux_stage_4[91] <= mux_stage_5[91]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[92] <= 0; else if(sel[4] == 1'b1) mux_stage_4[92] <= mux_stage_5[108]; else mux_stage_4[92] <= mux_stage_5[92]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[93] <= 0; else if(sel[4] == 1'b1) mux_stage_4[93] <= mux_stage_5[109]; else mux_stage_4[93] <= mux_stage_5[93]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[94] <= 0; else if(sel[4] == 1'b1) mux_stage_4[94] <= mux_stage_5[110]; else mux_stage_4[94] <= mux_stage_5[94]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[95] <= 0; else if(sel[4] == 1'b1) mux_stage_4[95] <= mux_stage_5[111]; else mux_stage_4[95] <= mux_stage_5[95]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[96] <= 0; else if(sel[4] == 1'b1) mux_stage_4[96] <= mux_stage_5[112]; else mux_stage_4[96] <= mux_stage_5[96]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[97] <= 0; else if(sel[4] == 1'b1) mux_stage_4[97] <= mux_stage_5[113]; else mux_stage_4[97] <= mux_stage_5[97]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[98] <= 0; else if(sel[4] == 1'b1) mux_stage_4[98] <= mux_stage_5[114]; else mux_stage_4[98] <= mux_stage_5[98]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[99] <= 0; else if(sel[4] == 1'b1) mux_stage_4[99] <= mux_stage_5[115]; else mux_stage_4[99] <= mux_stage_5[99]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[100] <= 0; else if(sel[4] == 1'b1) mux_stage_4[100] <= mux_stage_5[116]; else mux_stage_4[100] <= mux_stage_5[100]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[101] <= 0; else if(sel[4] == 1'b1) mux_stage_4[101] <= mux_stage_5[117]; else mux_stage_4[101] <= mux_stage_5[101]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[102] <= 0; else if(sel[4] == 1'b1) mux_stage_4[102] <= mux_stage_5[118]; else mux_stage_4[102] <= mux_stage_5[102]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[103] <= 0; else if(sel[4] == 1'b1) mux_stage_4[103] <= mux_stage_5[119]; else mux_stage_4[103] <= mux_stage_5[103]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[104] <= 0; else if(sel[4] == 1'b1) mux_stage_4[104] <= mux_stage_5[120]; else mux_stage_4[104] <= mux_stage_5[104]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[105] <= 0; else if(sel[4] == 1'b1) mux_stage_4[105] <= mux_stage_5[121]; else mux_stage_4[105] <= mux_stage_5[105]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[106] <= 0; else if(sel[4] == 1'b1) mux_stage_4[106] <= mux_stage_5[122]; else mux_stage_4[106] <= mux_stage_5[106]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[107] <= 0; else if(sel[4] == 1'b1) mux_stage_4[107] <= mux_stage_5[123]; else mux_stage_4[107] <= mux_stage_5[107]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[108] <= 0; else if(sel[4] == 1'b1) mux_stage_4[108] <= mux_stage_5[124]; else mux_stage_4[108] <= mux_stage_5[108]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[109] <= 0; else if(sel[4] == 1'b1) mux_stage_4[109] <= mux_stage_5[125]; else mux_stage_4[109] <= mux_stage_5[109]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[110] <= 0; else if(sel[4] == 1'b1) mux_stage_4[110] <= mux_stage_5[126]; else mux_stage_4[110] <= mux_stage_5[110]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[111] <= 0; else if(sel[4] == 1'b1) mux_stage_4[111] <= mux_stage_5[127]; else mux_stage_4[111] <= mux_stage_5[111]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[112] <= 0; else if(sel[4] == 1'b1) mux_stage_4[112] <= mux_stage_5[128]; else mux_stage_4[112] <= mux_stage_5[112]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[113] <= 0; else if(sel[4] == 1'b1) mux_stage_4[113] <= mux_stage_5[129]; else mux_stage_4[113] <= mux_stage_5[113]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[114] <= 0; else if(sel[4] == 1'b1) mux_stage_4[114] <= mux_stage_5[130]; else mux_stage_4[114] <= mux_stage_5[114]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[115] <= 0; else if(sel[4] == 1'b1) mux_stage_4[115] <= mux_stage_5[131]; else mux_stage_4[115] <= mux_stage_5[115]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[116] <= 0; else if(sel[4] == 1'b1) mux_stage_4[116] <= mux_stage_5[132]; else mux_stage_4[116] <= mux_stage_5[116]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[117] <= 0; else if(sel[4] == 1'b1) mux_stage_4[117] <= mux_stage_5[133]; else mux_stage_4[117] <= mux_stage_5[117]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[118] <= 0; else if(sel[4] == 1'b1) mux_stage_4[118] <= mux_stage_5[134]; else mux_stage_4[118] <= mux_stage_5[118]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[119] <= 0; else if(sel[4] == 1'b1) mux_stage_4[119] <= mux_stage_5[135]; else mux_stage_4[119] <= mux_stage_5[119]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[120] <= 0; else if(sel[4] == 1'b1) mux_stage_4[120] <= mux_stage_5[136]; else mux_stage_4[120] <= mux_stage_5[120]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[121] <= 0; else if(sel[4] == 1'b1) mux_stage_4[121] <= mux_stage_5[137]; else mux_stage_4[121] <= mux_stage_5[121]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[122] <= 0; else if(sel[4] == 1'b1) mux_stage_4[122] <= mux_stage_5[138]; else mux_stage_4[122] <= mux_stage_5[122]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[123] <= 0; else if(sel[4] == 1'b1) mux_stage_4[123] <= mux_stage_5[139]; else mux_stage_4[123] <= mux_stage_5[123]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[124] <= 0; else if(sel[4] == 1'b1) mux_stage_4[124] <= mux_stage_5[140]; else mux_stage_4[124] <= mux_stage_5[124]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[125] <= 0; else if(sel[4] == 1'b1) mux_stage_4[125] <= mux_stage_5[141]; else mux_stage_4[125] <= mux_stage_5[125]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[126] <= 0; else if(sel[4] == 1'b1) mux_stage_4[126] <= mux_stage_5[142]; else mux_stage_4[126] <= mux_stage_5[126]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[127] <= 0; else if(sel[4] == 1'b1) mux_stage_4[127] <= mux_stage_5[143]; else mux_stage_4[127] <= mux_stage_5[127]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[128] <= 0; else if(sel[4] == 1'b1) mux_stage_4[128] <= mux_stage_5[144]; else mux_stage_4[128] <= mux_stage_5[128]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[129] <= 0; else if(sel[4] == 1'b1) mux_stage_4[129] <= mux_stage_5[145]; else mux_stage_4[129] <= mux_stage_5[129]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[130] <= 0; else if(sel[4] == 1'b1) mux_stage_4[130] <= mux_stage_5[146]; else mux_stage_4[130] <= mux_stage_5[130]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[131] <= 0; else if(sel[4] == 1'b1) mux_stage_4[131] <= mux_stage_5[147]; else mux_stage_4[131] <= mux_stage_5[131]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[132] <= 0; else if(sel[4] == 1'b1) mux_stage_4[132] <= mux_stage_5[148]; else mux_stage_4[132] <= mux_stage_5[132]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[133] <= 0; else if(sel[4] == 1'b1) mux_stage_4[133] <= mux_stage_5[149]; else mux_stage_4[133] <= mux_stage_5[133]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[134] <= 0; else if(sel[4] == 1'b1) mux_stage_4[134] <= mux_stage_5[150]; else mux_stage_4[134] <= mux_stage_5[134]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[135] <= 0; else if(sel[4] == 1'b1) mux_stage_4[135] <= mux_stage_5[151]; else mux_stage_4[135] <= mux_stage_5[135]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[136] <= 0; else if(sel[4] == 1'b1) mux_stage_4[136] <= mux_stage_5[152]; else mux_stage_4[136] <= mux_stage_5[136]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[137] <= 0; else if(sel[4] == 1'b1) mux_stage_4[137] <= mux_stage_5[153]; else mux_stage_4[137] <= mux_stage_5[137]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[138] <= 0; else if(sel[4] == 1'b1) mux_stage_4[138] <= mux_stage_5[154]; else mux_stage_4[138] <= mux_stage_5[138]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[139] <= 0; else if(sel[4] == 1'b1) mux_stage_4[139] <= mux_stage_5[155]; else mux_stage_4[139] <= mux_stage_5[139]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[140] <= 0; else if(sel[4] == 1'b1) mux_stage_4[140] <= mux_stage_5[156]; else mux_stage_4[140] <= mux_stage_5[140]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[141] <= 0; else if(sel[4] == 1'b1) mux_stage_4[141] <= mux_stage_5[157]; else mux_stage_4[141] <= mux_stage_5[141]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[142] <= 0; else if(sel[4] == 1'b1) mux_stage_4[142] <= mux_stage_5[158]; else mux_stage_4[142] <= mux_stage_5[142]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[143] <= 0; else if(sel[4] == 1'b1) mux_stage_4[143] <= mux_stage_5[159]; else mux_stage_4[143] <= mux_stage_5[143]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[144] <= 0; else if(sel[4] == 1'b1) mux_stage_4[144] <= mux_stage_5[160]; else mux_stage_4[144] <= mux_stage_5[144]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[145] <= 0; else if(sel[4] == 1'b1) mux_stage_4[145] <= mux_stage_5[161]; else mux_stage_4[145] <= mux_stage_5[145]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[146] <= 0; else if(sel[4] == 1'b1) mux_stage_4[146] <= mux_stage_5[162]; else mux_stage_4[146] <= mux_stage_5[146]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[147] <= 0; else if(sel[4] == 1'b1) mux_stage_4[147] <= mux_stage_5[163]; else mux_stage_4[147] <= mux_stage_5[147]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[148] <= 0; else if(sel[4] == 1'b1) mux_stage_4[148] <= mux_stage_5[164]; else mux_stage_4[148] <= mux_stage_5[148]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[149] <= 0; else if(sel[4] == 1'b1) mux_stage_4[149] <= mux_stage_5[165]; else mux_stage_4[149] <= mux_stage_5[149]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[150] <= 0; else if(sel[4] == 1'b1) mux_stage_4[150] <= mux_stage_5[166]; else mux_stage_4[150] <= mux_stage_5[150]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[151] <= 0; else if(sel[4] == 1'b1) mux_stage_4[151] <= mux_stage_5[167]; else mux_stage_4[151] <= mux_stage_5[151]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[152] <= 0; else if(sel[4] == 1'b1) mux_stage_4[152] <= mux_stage_5[168]; else mux_stage_4[152] <= mux_stage_5[152]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[153] <= 0; else if(sel[4] == 1'b1) mux_stage_4[153] <= mux_stage_5[169]; else mux_stage_4[153] <= mux_stage_5[153]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[154] <= 0; else if(sel[4] == 1'b1) mux_stage_4[154] <= mux_stage_5[170]; else mux_stage_4[154] <= mux_stage_5[154]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[155] <= 0; else if(sel[4] == 1'b1) mux_stage_4[155] <= mux_stage_5[171]; else mux_stage_4[155] <= mux_stage_5[155]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[156] <= 0; else if(sel[4] == 1'b1) mux_stage_4[156] <= mux_stage_5[172]; else mux_stage_4[156] <= mux_stage_5[156]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[157] <= 0; else if(sel[4] == 1'b1) mux_stage_4[157] <= mux_stage_5[173]; else mux_stage_4[157] <= mux_stage_5[157]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[158] <= 0; else if(sel[4] == 1'b1) mux_stage_4[158] <= mux_stage_5[174]; else mux_stage_4[158] <= mux_stage_5[158]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[159] <= 0; else if(sel[4] == 1'b1) mux_stage_4[159] <= mux_stage_5[175]; else mux_stage_4[159] <= mux_stage_5[159]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[160] <= 0; else if(sel[4] == 1'b1) mux_stage_4[160] <= mux_stage_5[176]; else mux_stage_4[160] <= mux_stage_5[160]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[161] <= 0; else if(sel[4] == 1'b1) mux_stage_4[161] <= mux_stage_5[177]; else mux_stage_4[161] <= mux_stage_5[161]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[162] <= 0; else if(sel[4] == 1'b1) mux_stage_4[162] <= mux_stage_5[178]; else mux_stage_4[162] <= mux_stage_5[162]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[163] <= 0; else if(sel[4] == 1'b1) mux_stage_4[163] <= mux_stage_5[179]; else mux_stage_4[163] <= mux_stage_5[163]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[164] <= 0; else if(sel[4] == 1'b1) mux_stage_4[164] <= mux_stage_5[180]; else mux_stage_4[164] <= mux_stage_5[164]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[165] <= 0; else if(sel[4] == 1'b1) mux_stage_4[165] <= mux_stage_5[181]; else mux_stage_4[165] <= mux_stage_5[165]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[166] <= 0; else if(sel[4] == 1'b1) mux_stage_4[166] <= mux_stage_5[182]; else mux_stage_4[166] <= mux_stage_5[166]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[167] <= 0; else if(sel[4] == 1'b1) mux_stage_4[167] <= mux_stage_5[183]; else mux_stage_4[167] <= mux_stage_5[167]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[168] <= 0; else if(sel[4] == 1'b1) mux_stage_4[168] <= mux_stage_5[184]; else mux_stage_4[168] <= mux_stage_5[168]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[169] <= 0; else if(sel[4] == 1'b1) mux_stage_4[169] <= mux_stage_5[185]; else mux_stage_4[169] <= mux_stage_5[169]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[170] <= 0; else if(sel[4] == 1'b1) mux_stage_4[170] <= mux_stage_5[186]; else mux_stage_4[170] <= mux_stage_5[170]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[171] <= 0; else if(sel[4] == 1'b1) mux_stage_4[171] <= mux_stage_5[187]; else mux_stage_4[171] <= mux_stage_5[171]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[172] <= 0; else if(sel[4] == 1'b1) mux_stage_4[172] <= mux_stage_5[188]; else mux_stage_4[172] <= mux_stage_5[172]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[173] <= 0; else if(sel[4] == 1'b1) mux_stage_4[173] <= mux_stage_5[189]; else mux_stage_4[173] <= mux_stage_5[173]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[174] <= 0; else if(sel[4] == 1'b1) mux_stage_4[174] <= mux_stage_5[190]; else mux_stage_4[174] <= mux_stage_5[174]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[175] <= 0; else if(sel[4] == 1'b1) mux_stage_4[175] <= mux_stage_5[191]; else mux_stage_4[175] <= mux_stage_5[175]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[176] <= 0; else if(sel[4] == 1'b1) mux_stage_4[176] <= mux_stage_5[192]; else mux_stage_4[176] <= mux_stage_5[176]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[177] <= 0; else if(sel[4] == 1'b1) mux_stage_4[177] <= mux_stage_5[193]; else mux_stage_4[177] <= mux_stage_5[177]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[178] <= 0; else if(sel[4] == 1'b1) mux_stage_4[178] <= mux_stage_5[194]; else mux_stage_4[178] <= mux_stage_5[178]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[179] <= 0; else if(sel[4] == 1'b1) mux_stage_4[179] <= mux_stage_5[195]; else mux_stage_4[179] <= mux_stage_5[179]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[180] <= 0; else if(sel[4] == 1'b1) mux_stage_4[180] <= mux_stage_5[196]; else mux_stage_4[180] <= mux_stage_5[180]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[181] <= 0; else if(sel[4] == 1'b1) mux_stage_4[181] <= mux_stage_5[197]; else mux_stage_4[181] <= mux_stage_5[181]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[182] <= 0; else if(sel[4] == 1'b1) mux_stage_4[182] <= mux_stage_5[198]; else mux_stage_4[182] <= mux_stage_5[182]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[183] <= 0; else if(sel[4] == 1'b1) mux_stage_4[183] <= mux_stage_5[199]; else mux_stage_4[183] <= mux_stage_5[183]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[184] <= 0; else if(sel[4] == 1'b1) mux_stage_4[184] <= mux_stage_5[200]; else mux_stage_4[184] <= mux_stage_5[184]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[185] <= 0; else if(sel[4] == 1'b1) mux_stage_4[185] <= mux_stage_5[201]; else mux_stage_4[185] <= mux_stage_5[185]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[186] <= 0; else if(sel[4] == 1'b1) mux_stage_4[186] <= mux_stage_5[202]; else mux_stage_4[186] <= mux_stage_5[186]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[187] <= 0; else if(sel[4] == 1'b1) mux_stage_4[187] <= mux_stage_5[203]; else mux_stage_4[187] <= mux_stage_5[187]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[188] <= 0; else if(sel[4] == 1'b1) mux_stage_4[188] <= mux_stage_5[204]; else mux_stage_4[188] <= mux_stage_5[188]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[189] <= 0; else if(sel[4] == 1'b1) mux_stage_4[189] <= mux_stage_5[205]; else mux_stage_4[189] <= mux_stage_5[189]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[190] <= 0; else if(sel[4] == 1'b1) mux_stage_4[190] <= mux_stage_5[206]; else mux_stage_4[190] <= mux_stage_5[190]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[191] <= 0; else if(sel[4] == 1'b1) mux_stage_4[191] <= mux_stage_5[207]; else mux_stage_4[191] <= mux_stage_5[191]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[192] <= 0; else if(sel[4] == 1'b1) mux_stage_4[192] <= mux_stage_5[208]; else mux_stage_4[192] <= mux_stage_5[192]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[193] <= 0; else if(sel[4] == 1'b1) mux_stage_4[193] <= mux_stage_5[209]; else mux_stage_4[193] <= mux_stage_5[193]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[194] <= 0; else if(sel[4] == 1'b1) mux_stage_4[194] <= mux_stage_5[210]; else mux_stage_4[194] <= mux_stage_5[194]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[195] <= 0; else if(sel[4] == 1'b1) mux_stage_4[195] <= mux_stage_5[211]; else mux_stage_4[195] <= mux_stage_5[195]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[196] <= 0; else if(sel[4] == 1'b1) mux_stage_4[196] <= mux_stage_5[212]; else mux_stage_4[196] <= mux_stage_5[196]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[197] <= 0; else if(sel[4] == 1'b1) mux_stage_4[197] <= mux_stage_5[213]; else mux_stage_4[197] <= mux_stage_5[197]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[198] <= 0; else if(sel[4] == 1'b1) mux_stage_4[198] <= mux_stage_5[214]; else mux_stage_4[198] <= mux_stage_5[198]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[199] <= 0; else if(sel[4] == 1'b1) mux_stage_4[199] <= mux_stage_5[215]; else mux_stage_4[199] <= mux_stage_5[199]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[200] <= 0; else if(sel[4] == 1'b1) mux_stage_4[200] <= mux_stage_5[216]; else mux_stage_4[200] <= mux_stage_5[200]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[201] <= 0; else if(sel[4] == 1'b1) mux_stage_4[201] <= mux_stage_5[217]; else mux_stage_4[201] <= mux_stage_5[201]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[202] <= 0; else if(sel[4] == 1'b1) mux_stage_4[202] <= mux_stage_5[218]; else mux_stage_4[202] <= mux_stage_5[202]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[203] <= 0; else if(sel[4] == 1'b1) mux_stage_4[203] <= mux_stage_5[219]; else mux_stage_4[203] <= mux_stage_5[203]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[204] <= 0; else if(sel[4] == 1'b1) mux_stage_4[204] <= mux_stage_5[220]; else mux_stage_4[204] <= mux_stage_5[204]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[205] <= 0; else if(sel[4] == 1'b1) mux_stage_4[205] <= mux_stage_5[221]; else mux_stage_4[205] <= mux_stage_5[205]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[206] <= 0; else if(sel[4] == 1'b1) mux_stage_4[206] <= mux_stage_5[222]; else mux_stage_4[206] <= mux_stage_5[206]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[207] <= 0; else if(sel[4] == 1'b1) mux_stage_4[207] <= sw_in[223]; else mux_stage_4[207] <= mux_stage_5[207]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[208] <= 0; else if(sel[4] == 1'b1) mux_stage_4[208] <= sw_in[224]; else mux_stage_4[208] <= mux_stage_5[208]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[209] <= 0; else if(sel[4] == 1'b1) mux_stage_4[209] <= sw_in[225]; else mux_stage_4[209] <= mux_stage_5[209]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[210] <= 0; else if(sel[4] == 1'b1) mux_stage_4[210] <= sw_in[226]; else mux_stage_4[210] <= mux_stage_5[210]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[211] <= 0; else if(sel[4] == 1'b1) mux_stage_4[211] <= sw_in[227]; else mux_stage_4[211] <= mux_stage_5[211]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[212] <= 0; else if(sel[4] == 1'b1) mux_stage_4[212] <= sw_in[228]; else mux_stage_4[212] <= mux_stage_5[212]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[213] <= 0; else if(sel[4] == 1'b1) mux_stage_4[213] <= sw_in[229]; else mux_stage_4[213] <= mux_stage_5[213]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[214] <= 0; else if(sel[4] == 1'b1) mux_stage_4[214] <= sw_in[230]; else mux_stage_4[214] <= mux_stage_5[214]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[215] <= 0; else if(sel[4] == 1'b1) mux_stage_4[215] <= sw_in[231]; else mux_stage_4[215] <= mux_stage_5[215]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[216] <= 0; else if(sel[4] == 1'b1) mux_stage_4[216] <= sw_in[232]; else mux_stage_4[216] <= mux_stage_5[216]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[217] <= 0; else if(sel[4] == 1'b1) mux_stage_4[217] <= sw_in[233]; else mux_stage_4[217] <= mux_stage_5[217]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[218] <= 0; else if(sel[4] == 1'b1) mux_stage_4[218] <= sw_in[234]; else mux_stage_4[218] <= mux_stage_5[218]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[219] <= 0; else if(sel[4] == 1'b1) mux_stage_4[219] <= sw_in[235]; else mux_stage_4[219] <= mux_stage_5[219]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[220] <= 0; else if(sel[4] == 1'b1) mux_stage_4[220] <= sw_in[236]; else mux_stage_4[220] <= mux_stage_5[220]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[221] <= 0; else if(sel[4] == 1'b1) mux_stage_4[221] <= sw_in[237]; else mux_stage_4[221] <= mux_stage_5[221]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[222] <= 0; else if(sel[4] == 1'b1) mux_stage_4[222] <= sw_in[238]; else mux_stage_4[222] <= mux_stage_5[222]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[223] <= 0; else if(sel[4] == 1'b1) mux_stage_4[223] <= sw_in[239]; else mux_stage_4[223] <= sw_in[223]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[224] <= 0; else if(sel[4] == 1'b1) mux_stage_4[224] <= sw_in[240]; else mux_stage_4[224] <= sw_in[224]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[225] <= 0; else if(sel[4] == 1'b1) mux_stage_4[225] <= sw_in[241]; else mux_stage_4[225] <= sw_in[225]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[226] <= 0; else if(sel[4] == 1'b1) mux_stage_4[226] <= sw_in[242]; else mux_stage_4[226] <= sw_in[226]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[227] <= 0; else if(sel[4] == 1'b1) mux_stage_4[227] <= sw_in[243]; else mux_stage_4[227] <= sw_in[227]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[228] <= 0; else if(sel[4] == 1'b1) mux_stage_4[228] <= sw_in[244]; else mux_stage_4[228] <= sw_in[228]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[229] <= 0; else if(sel[4] == 1'b1) mux_stage_4[229] <= sw_in[245]; else mux_stage_4[229] <= sw_in[229]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[230] <= 0; else if(sel[4] == 1'b1) mux_stage_4[230] <= sw_in[246]; else mux_stage_4[230] <= sw_in[230]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[231] <= 0; else if(sel[4] == 1'b1) mux_stage_4[231] <= sw_in[247]; else mux_stage_4[231] <= sw_in[231]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[232] <= 0; else if(sel[4] == 1'b1) mux_stage_4[232] <= sw_in[248]; else mux_stage_4[232] <= sw_in[232]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[233] <= 0; else if(sel[4] == 1'b1) mux_stage_4[233] <= sw_in[249]; else mux_stage_4[233] <= sw_in[233]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[234] <= 0; else if(sel[4] == 1'b1) mux_stage_4[234] <= sw_in[250]; else mux_stage_4[234] <= sw_in[234]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[235] <= 0; else if(sel[4] == 1'b1) mux_stage_4[235] <= sw_in[251]; else mux_stage_4[235] <= sw_in[235]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[236] <= 0; else if(sel[4] == 1'b1) mux_stage_4[236] <= sw_in[252]; else mux_stage_4[236] <= sw_in[236]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[237] <= 0; else if(sel[4] == 1'b1) mux_stage_4[237] <= sw_in[253]; else mux_stage_4[237] <= sw_in[237]; end
	always @(posedge sys_clk) begin if(!rstn) mux_stage_4[238] <= 0; else if(sel[4] == 1'b1) mux_stage_4[238] <= sw_in[254]; else mux_stage_4[238] <= sw_in[238]; end

	reg sw_in_239_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_239_reg0 <= 0; else sw_in_239_reg0 <= sw_in[239]; end
	reg sw_in_240_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_240_reg0 <= 0; else sw_in_240_reg0 <= sw_in[240]; end
	reg sw_in_241_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_241_reg0 <= 0; else sw_in_241_reg0 <= sw_in[241]; end
	reg sw_in_242_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_242_reg0 <= 0; else sw_in_242_reg0 <= sw_in[242]; end
	reg sw_in_243_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_243_reg0 <= 0; else sw_in_243_reg0 <= sw_in[243]; end
	reg sw_in_244_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_244_reg0 <= 0; else sw_in_244_reg0 <= sw_in[244]; end
	reg sw_in_245_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_245_reg0 <= 0; else sw_in_245_reg0 <= sw_in[245]; end
	reg sw_in_246_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_246_reg0 <= 0; else sw_in_246_reg0 <= sw_in[246]; end
	reg sw_in_247_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_247_reg0 <= 0; else sw_in_247_reg0 <= sw_in[247]; end
	reg sw_in_248_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_248_reg0 <= 0; else sw_in_248_reg0 <= sw_in[248]; end
	reg sw_in_249_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_249_reg0 <= 0; else sw_in_249_reg0 <= sw_in[249]; end
	reg sw_in_250_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_250_reg0 <= 0; else sw_in_250_reg0 <= sw_in[250]; end
	reg sw_in_251_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_251_reg0 <= 0; else sw_in_251_reg0 <= sw_in[251]; end
	reg sw_in_252_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_252_reg0 <= 0; else sw_in_252_reg0 <= sw_in[252]; end
	reg sw_in_253_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_253_reg0 <= 0; else sw_in_253_reg0 <= sw_in[253]; end
	reg sw_in_254_reg0; 	always @(posedge sys_clk) begin if(!rstn) sw_in_254_reg0 <= 0; else sw_in_254_reg0 <= sw_in[254]; end

	reg sel_3_reg0;
	always @(posedge sys_clk) begin if(!rstn) sel_3_reg0 <= 0; else sel_3_reg0 <= sel[3]; end	

	// Multiplexer Stage 3
	wire [246:0] mux_stage_3;
	assign mux_stage_3[0] = (sel_3_reg0 == 1'b1) ? mux_stage_4[8] : mux_stage_4[0];
	assign mux_stage_3[1] = (sel_3_reg0 == 1'b1) ? mux_stage_4[9] : mux_stage_4[1];
	assign mux_stage_3[2] = (sel_3_reg0 == 1'b1) ? mux_stage_4[10] : mux_stage_4[2];
	assign mux_stage_3[3] = (sel_3_reg0 == 1'b1) ? mux_stage_4[11] : mux_stage_4[3];
	assign mux_stage_3[4] = (sel_3_reg0 == 1'b1) ? mux_stage_4[12] : mux_stage_4[4];
	assign mux_stage_3[5] = (sel_3_reg0 == 1'b1) ? mux_stage_4[13] : mux_stage_4[5];
	assign mux_stage_3[6] = (sel_3_reg0 == 1'b1) ? mux_stage_4[14] : mux_stage_4[6];
	assign mux_stage_3[7] = (sel_3_reg0 == 1'b1) ? mux_stage_4[15] : mux_stage_4[7];
	assign mux_stage_3[8] = (sel_3_reg0 == 1'b1) ? mux_stage_4[16] : mux_stage_4[8];
	assign mux_stage_3[9] = (sel_3_reg0 == 1'b1) ? mux_stage_4[17] : mux_stage_4[9];
	assign mux_stage_3[10] = (sel_3_reg0 == 1'b1) ? mux_stage_4[18] : mux_stage_4[10];
	assign mux_stage_3[11] = (sel_3_reg0 == 1'b1) ? mux_stage_4[19] : mux_stage_4[11];
	assign mux_stage_3[12] = (sel_3_reg0 == 1'b1) ? mux_stage_4[20] : mux_stage_4[12];
	assign mux_stage_3[13] = (sel_3_reg0 == 1'b1) ? mux_stage_4[21] : mux_stage_4[13];
	assign mux_stage_3[14] = (sel_3_reg0 == 1'b1) ? mux_stage_4[22] : mux_stage_4[14];
	assign mux_stage_3[15] = (sel_3_reg0 == 1'b1) ? mux_stage_4[23] : mux_stage_4[15];
	assign mux_stage_3[16] = (sel_3_reg0 == 1'b1) ? mux_stage_4[24] : mux_stage_4[16];
	assign mux_stage_3[17] = (sel_3_reg0 == 1'b1) ? mux_stage_4[25] : mux_stage_4[17];
	assign mux_stage_3[18] = (sel_3_reg0 == 1'b1) ? mux_stage_4[26] : mux_stage_4[18];
	assign mux_stage_3[19] = (sel_3_reg0 == 1'b1) ? mux_stage_4[27] : mux_stage_4[19];
	assign mux_stage_3[20] = (sel_3_reg0 == 1'b1) ? mux_stage_4[28] : mux_stage_4[20];
	assign mux_stage_3[21] = (sel_3_reg0 == 1'b1) ? mux_stage_4[29] : mux_stage_4[21];
	assign mux_stage_3[22] = (sel_3_reg0 == 1'b1) ? mux_stage_4[30] : mux_stage_4[22];
	assign mux_stage_3[23] = (sel_3_reg0 == 1'b1) ? mux_stage_4[31] : mux_stage_4[23];
	assign mux_stage_3[24] = (sel_3_reg0 == 1'b1) ? mux_stage_4[32] : mux_stage_4[24];
	assign mux_stage_3[25] = (sel_3_reg0 == 1'b1) ? mux_stage_4[33] : mux_stage_4[25];
	assign mux_stage_3[26] = (sel_3_reg0 == 1'b1) ? mux_stage_4[34] : mux_stage_4[26];
	assign mux_stage_3[27] = (sel_3_reg0 == 1'b1) ? mux_stage_4[35] : mux_stage_4[27];
	assign mux_stage_3[28] = (sel_3_reg0 == 1'b1) ? mux_stage_4[36] : mux_stage_4[28];
	assign mux_stage_3[29] = (sel_3_reg0 == 1'b1) ? mux_stage_4[37] : mux_stage_4[29];
	assign mux_stage_3[30] = (sel_3_reg0 == 1'b1) ? mux_stage_4[38] : mux_stage_4[30];
	assign mux_stage_3[31] = (sel_3_reg0 == 1'b1) ? mux_stage_4[39] : mux_stage_4[31];
	assign mux_stage_3[32] = (sel_3_reg0 == 1'b1) ? mux_stage_4[40] : mux_stage_4[32];
	assign mux_stage_3[33] = (sel_3_reg0 == 1'b1) ? mux_stage_4[41] : mux_stage_4[33];
	assign mux_stage_3[34] = (sel_3_reg0 == 1'b1) ? mux_stage_4[42] : mux_stage_4[34];
	assign mux_stage_3[35] = (sel_3_reg0 == 1'b1) ? mux_stage_4[43] : mux_stage_4[35];
	assign mux_stage_3[36] = (sel_3_reg0 == 1'b1) ? mux_stage_4[44] : mux_stage_4[36];
	assign mux_stage_3[37] = (sel_3_reg0 == 1'b1) ? mux_stage_4[45] : mux_stage_4[37];
	assign mux_stage_3[38] = (sel_3_reg0 == 1'b1) ? mux_stage_4[46] : mux_stage_4[38];
	assign mux_stage_3[39] = (sel_3_reg0 == 1'b1) ? mux_stage_4[47] : mux_stage_4[39];
	assign mux_stage_3[40] = (sel_3_reg0 == 1'b1) ? mux_stage_4[48] : mux_stage_4[40];
	assign mux_stage_3[41] = (sel_3_reg0 == 1'b1) ? mux_stage_4[49] : mux_stage_4[41];
	assign mux_stage_3[42] = (sel_3_reg0 == 1'b1) ? mux_stage_4[50] : mux_stage_4[42];
	assign mux_stage_3[43] = (sel_3_reg0 == 1'b1) ? mux_stage_4[51] : mux_stage_4[43];
	assign mux_stage_3[44] = (sel_3_reg0 == 1'b1) ? mux_stage_4[52] : mux_stage_4[44];
	assign mux_stage_3[45] = (sel_3_reg0 == 1'b1) ? mux_stage_4[53] : mux_stage_4[45];
	assign mux_stage_3[46] = (sel_3_reg0 == 1'b1) ? mux_stage_4[54] : mux_stage_4[46];
	assign mux_stage_3[47] = (sel_3_reg0 == 1'b1) ? mux_stage_4[55] : mux_stage_4[47];
	assign mux_stage_3[48] = (sel_3_reg0 == 1'b1) ? mux_stage_4[56] : mux_stage_4[48];
	assign mux_stage_3[49] = (sel_3_reg0 == 1'b1) ? mux_stage_4[57] : mux_stage_4[49];
	assign mux_stage_3[50] = (sel_3_reg0 == 1'b1) ? mux_stage_4[58] : mux_stage_4[50];
	assign mux_stage_3[51] = (sel_3_reg0 == 1'b1) ? mux_stage_4[59] : mux_stage_4[51];
	assign mux_stage_3[52] = (sel_3_reg0 == 1'b1) ? mux_stage_4[60] : mux_stage_4[52];
	assign mux_stage_3[53] = (sel_3_reg0 == 1'b1) ? mux_stage_4[61] : mux_stage_4[53];
	assign mux_stage_3[54] = (sel_3_reg0 == 1'b1) ? mux_stage_4[62] : mux_stage_4[54];
	assign mux_stage_3[55] = (sel_3_reg0 == 1'b1) ? mux_stage_4[63] : mux_stage_4[55];
	assign mux_stage_3[56] = (sel_3_reg0 == 1'b1) ? mux_stage_4[64] : mux_stage_4[56];
	assign mux_stage_3[57] = (sel_3_reg0 == 1'b1) ? mux_stage_4[65] : mux_stage_4[57];
	assign mux_stage_3[58] = (sel_3_reg0 == 1'b1) ? mux_stage_4[66] : mux_stage_4[58];
	assign mux_stage_3[59] = (sel_3_reg0 == 1'b1) ? mux_stage_4[67] : mux_stage_4[59];
	assign mux_stage_3[60] = (sel_3_reg0 == 1'b1) ? mux_stage_4[68] : mux_stage_4[60];
	assign mux_stage_3[61] = (sel_3_reg0 == 1'b1) ? mux_stage_4[69] : mux_stage_4[61];
	assign mux_stage_3[62] = (sel_3_reg0 == 1'b1) ? mux_stage_4[70] : mux_stage_4[62];
	assign mux_stage_3[63] = (sel_3_reg0 == 1'b1) ? mux_stage_4[71] : mux_stage_4[63];
	assign mux_stage_3[64] = (sel_3_reg0 == 1'b1) ? mux_stage_4[72] : mux_stage_4[64];
	assign mux_stage_3[65] = (sel_3_reg0 == 1'b1) ? mux_stage_4[73] : mux_stage_4[65];
	assign mux_stage_3[66] = (sel_3_reg0 == 1'b1) ? mux_stage_4[74] : mux_stage_4[66];
	assign mux_stage_3[67] = (sel_3_reg0 == 1'b1) ? mux_stage_4[75] : mux_stage_4[67];
	assign mux_stage_3[68] = (sel_3_reg0 == 1'b1) ? mux_stage_4[76] : mux_stage_4[68];
	assign mux_stage_3[69] = (sel_3_reg0 == 1'b1) ? mux_stage_4[77] : mux_stage_4[69];
	assign mux_stage_3[70] = (sel_3_reg0 == 1'b1) ? mux_stage_4[78] : mux_stage_4[70];
	assign mux_stage_3[71] = (sel_3_reg0 == 1'b1) ? mux_stage_4[79] : mux_stage_4[71];
	assign mux_stage_3[72] = (sel_3_reg0 == 1'b1) ? mux_stage_4[80] : mux_stage_4[72];
	assign mux_stage_3[73] = (sel_3_reg0 == 1'b1) ? mux_stage_4[81] : mux_stage_4[73];
	assign mux_stage_3[74] = (sel_3_reg0 == 1'b1) ? mux_stage_4[82] : mux_stage_4[74];
	assign mux_stage_3[75] = (sel_3_reg0 == 1'b1) ? mux_stage_4[83] : mux_stage_4[75];
	assign mux_stage_3[76] = (sel_3_reg0 == 1'b1) ? mux_stage_4[84] : mux_stage_4[76];
	assign mux_stage_3[77] = (sel_3_reg0 == 1'b1) ? mux_stage_4[85] : mux_stage_4[77];
	assign mux_stage_3[78] = (sel_3_reg0 == 1'b1) ? mux_stage_4[86] : mux_stage_4[78];
	assign mux_stage_3[79] = (sel_3_reg0 == 1'b1) ? mux_stage_4[87] : mux_stage_4[79];
	assign mux_stage_3[80] = (sel_3_reg0 == 1'b1) ? mux_stage_4[88] : mux_stage_4[80];
	assign mux_stage_3[81] = (sel_3_reg0 == 1'b1) ? mux_stage_4[89] : mux_stage_4[81];
	assign mux_stage_3[82] = (sel_3_reg0 == 1'b1) ? mux_stage_4[90] : mux_stage_4[82];
	assign mux_stage_3[83] = (sel_3_reg0 == 1'b1) ? mux_stage_4[91] : mux_stage_4[83];
	assign mux_stage_3[84] = (sel_3_reg0 == 1'b1) ? mux_stage_4[92] : mux_stage_4[84];
	assign mux_stage_3[85] = (sel_3_reg0 == 1'b1) ? mux_stage_4[93] : mux_stage_4[85];
	assign mux_stage_3[86] = (sel_3_reg0 == 1'b1) ? mux_stage_4[94] : mux_stage_4[86];
	assign mux_stage_3[87] = (sel_3_reg0 == 1'b1) ? mux_stage_4[95] : mux_stage_4[87];
	assign mux_stage_3[88] = (sel_3_reg0 == 1'b1) ? mux_stage_4[96] : mux_stage_4[88];
	assign mux_stage_3[89] = (sel_3_reg0 == 1'b1) ? mux_stage_4[97] : mux_stage_4[89];
	assign mux_stage_3[90] = (sel_3_reg0 == 1'b1) ? mux_stage_4[98] : mux_stage_4[90];
	assign mux_stage_3[91] = (sel_3_reg0 == 1'b1) ? mux_stage_4[99] : mux_stage_4[91];
	assign mux_stage_3[92] = (sel_3_reg0 == 1'b1) ? mux_stage_4[100] : mux_stage_4[92];
	assign mux_stage_3[93] = (sel_3_reg0 == 1'b1) ? mux_stage_4[101] : mux_stage_4[93];
	assign mux_stage_3[94] = (sel_3_reg0 == 1'b1) ? mux_stage_4[102] : mux_stage_4[94];
	assign mux_stage_3[95] = (sel_3_reg0 == 1'b1) ? mux_stage_4[103] : mux_stage_4[95];
	assign mux_stage_3[96] = (sel_3_reg0 == 1'b1) ? mux_stage_4[104] : mux_stage_4[96];
	assign mux_stage_3[97] = (sel_3_reg0 == 1'b1) ? mux_stage_4[105] : mux_stage_4[97];
	assign mux_stage_3[98] = (sel_3_reg0 == 1'b1) ? mux_stage_4[106] : mux_stage_4[98];
	assign mux_stage_3[99] = (sel_3_reg0 == 1'b1) ? mux_stage_4[107] : mux_stage_4[99];
	assign mux_stage_3[100] = (sel_3_reg0 == 1'b1) ? mux_stage_4[108] : mux_stage_4[100];
	assign mux_stage_3[101] = (sel_3_reg0 == 1'b1) ? mux_stage_4[109] : mux_stage_4[101];
	assign mux_stage_3[102] = (sel_3_reg0 == 1'b1) ? mux_stage_4[110] : mux_stage_4[102];
	assign mux_stage_3[103] = (sel_3_reg0 == 1'b1) ? mux_stage_4[111] : mux_stage_4[103];
	assign mux_stage_3[104] = (sel_3_reg0 == 1'b1) ? mux_stage_4[112] : mux_stage_4[104];
	assign mux_stage_3[105] = (sel_3_reg0 == 1'b1) ? mux_stage_4[113] : mux_stage_4[105];
	assign mux_stage_3[106] = (sel_3_reg0 == 1'b1) ? mux_stage_4[114] : mux_stage_4[106];
	assign mux_stage_3[107] = (sel_3_reg0 == 1'b1) ? mux_stage_4[115] : mux_stage_4[107];
	assign mux_stage_3[108] = (sel_3_reg0 == 1'b1) ? mux_stage_4[116] : mux_stage_4[108];
	assign mux_stage_3[109] = (sel_3_reg0 == 1'b1) ? mux_stage_4[117] : mux_stage_4[109];
	assign mux_stage_3[110] = (sel_3_reg0 == 1'b1) ? mux_stage_4[118] : mux_stage_4[110];
	assign mux_stage_3[111] = (sel_3_reg0 == 1'b1) ? mux_stage_4[119] : mux_stage_4[111];
	assign mux_stage_3[112] = (sel_3_reg0 == 1'b1) ? mux_stage_4[120] : mux_stage_4[112];
	assign mux_stage_3[113] = (sel_3_reg0 == 1'b1) ? mux_stage_4[121] : mux_stage_4[113];
	assign mux_stage_3[114] = (sel_3_reg0 == 1'b1) ? mux_stage_4[122] : mux_stage_4[114];
	assign mux_stage_3[115] = (sel_3_reg0 == 1'b1) ? mux_stage_4[123] : mux_stage_4[115];
	assign mux_stage_3[116] = (sel_3_reg0 == 1'b1) ? mux_stage_4[124] : mux_stage_4[116];
	assign mux_stage_3[117] = (sel_3_reg0 == 1'b1) ? mux_stage_4[125] : mux_stage_4[117];
	assign mux_stage_3[118] = (sel_3_reg0 == 1'b1) ? mux_stage_4[126] : mux_stage_4[118];
	assign mux_stage_3[119] = (sel_3_reg0 == 1'b1) ? mux_stage_4[127] : mux_stage_4[119];
	assign mux_stage_3[120] = (sel_3_reg0 == 1'b1) ? mux_stage_4[128] : mux_stage_4[120];
	assign mux_stage_3[121] = (sel_3_reg0 == 1'b1) ? mux_stage_4[129] : mux_stage_4[121];
	assign mux_stage_3[122] = (sel_3_reg0 == 1'b1) ? mux_stage_4[130] : mux_stage_4[122];
	assign mux_stage_3[123] = (sel_3_reg0 == 1'b1) ? mux_stage_4[131] : mux_stage_4[123];
	assign mux_stage_3[124] = (sel_3_reg0 == 1'b1) ? mux_stage_4[132] : mux_stage_4[124];
	assign mux_stage_3[125] = (sel_3_reg0 == 1'b1) ? mux_stage_4[133] : mux_stage_4[125];
	assign mux_stage_3[126] = (sel_3_reg0 == 1'b1) ? mux_stage_4[134] : mux_stage_4[126];
	assign mux_stage_3[127] = (sel_3_reg0 == 1'b1) ? mux_stage_4[135] : mux_stage_4[127];
	assign mux_stage_3[128] = (sel_3_reg0 == 1'b1) ? mux_stage_4[136] : mux_stage_4[128];
	assign mux_stage_3[129] = (sel_3_reg0 == 1'b1) ? mux_stage_4[137] : mux_stage_4[129];
	assign mux_stage_3[130] = (sel_3_reg0 == 1'b1) ? mux_stage_4[138] : mux_stage_4[130];
	assign mux_stage_3[131] = (sel_3_reg0 == 1'b1) ? mux_stage_4[139] : mux_stage_4[131];
	assign mux_stage_3[132] = (sel_3_reg0 == 1'b1) ? mux_stage_4[140] : mux_stage_4[132];
	assign mux_stage_3[133] = (sel_3_reg0 == 1'b1) ? mux_stage_4[141] : mux_stage_4[133];
	assign mux_stage_3[134] = (sel_3_reg0 == 1'b1) ? mux_stage_4[142] : mux_stage_4[134];
	assign mux_stage_3[135] = (sel_3_reg0 == 1'b1) ? mux_stage_4[143] : mux_stage_4[135];
	assign mux_stage_3[136] = (sel_3_reg0 == 1'b1) ? mux_stage_4[144] : mux_stage_4[136];
	assign mux_stage_3[137] = (sel_3_reg0 == 1'b1) ? mux_stage_4[145] : mux_stage_4[137];
	assign mux_stage_3[138] = (sel_3_reg0 == 1'b1) ? mux_stage_4[146] : mux_stage_4[138];
	assign mux_stage_3[139] = (sel_3_reg0 == 1'b1) ? mux_stage_4[147] : mux_stage_4[139];
	assign mux_stage_3[140] = (sel_3_reg0 == 1'b1) ? mux_stage_4[148] : mux_stage_4[140];
	assign mux_stage_3[141] = (sel_3_reg0 == 1'b1) ? mux_stage_4[149] : mux_stage_4[141];
	assign mux_stage_3[142] = (sel_3_reg0 == 1'b1) ? mux_stage_4[150] : mux_stage_4[142];
	assign mux_stage_3[143] = (sel_3_reg0 == 1'b1) ? mux_stage_4[151] : mux_stage_4[143];
	assign mux_stage_3[144] = (sel_3_reg0 == 1'b1) ? mux_stage_4[152] : mux_stage_4[144];
	assign mux_stage_3[145] = (sel_3_reg0 == 1'b1) ? mux_stage_4[153] : mux_stage_4[145];
	assign mux_stage_3[146] = (sel_3_reg0 == 1'b1) ? mux_stage_4[154] : mux_stage_4[146];
	assign mux_stage_3[147] = (sel_3_reg0 == 1'b1) ? mux_stage_4[155] : mux_stage_4[147];
	assign mux_stage_3[148] = (sel_3_reg0 == 1'b1) ? mux_stage_4[156] : mux_stage_4[148];
	assign mux_stage_3[149] = (sel_3_reg0 == 1'b1) ? mux_stage_4[157] : mux_stage_4[149];
	assign mux_stage_3[150] = (sel_3_reg0 == 1'b1) ? mux_stage_4[158] : mux_stage_4[150];
	assign mux_stage_3[151] = (sel_3_reg0 == 1'b1) ? mux_stage_4[159] : mux_stage_4[151];
	assign mux_stage_3[152] = (sel_3_reg0 == 1'b1) ? mux_stage_4[160] : mux_stage_4[152];
	assign mux_stage_3[153] = (sel_3_reg0 == 1'b1) ? mux_stage_4[161] : mux_stage_4[153];
	assign mux_stage_3[154] = (sel_3_reg0 == 1'b1) ? mux_stage_4[162] : mux_stage_4[154];
	assign mux_stage_3[155] = (sel_3_reg0 == 1'b1) ? mux_stage_4[163] : mux_stage_4[155];
	assign mux_stage_3[156] = (sel_3_reg0 == 1'b1) ? mux_stage_4[164] : mux_stage_4[156];
	assign mux_stage_3[157] = (sel_3_reg0 == 1'b1) ? mux_stage_4[165] : mux_stage_4[157];
	assign mux_stage_3[158] = (sel_3_reg0 == 1'b1) ? mux_stage_4[166] : mux_stage_4[158];
	assign mux_stage_3[159] = (sel_3_reg0 == 1'b1) ? mux_stage_4[167] : mux_stage_4[159];
	assign mux_stage_3[160] = (sel_3_reg0 == 1'b1) ? mux_stage_4[168] : mux_stage_4[160];
	assign mux_stage_3[161] = (sel_3_reg0 == 1'b1) ? mux_stage_4[169] : mux_stage_4[161];
	assign mux_stage_3[162] = (sel_3_reg0 == 1'b1) ? mux_stage_4[170] : mux_stage_4[162];
	assign mux_stage_3[163] = (sel_3_reg0 == 1'b1) ? mux_stage_4[171] : mux_stage_4[163];
	assign mux_stage_3[164] = (sel_3_reg0 == 1'b1) ? mux_stage_4[172] : mux_stage_4[164];
	assign mux_stage_3[165] = (sel_3_reg0 == 1'b1) ? mux_stage_4[173] : mux_stage_4[165];
	assign mux_stage_3[166] = (sel_3_reg0 == 1'b1) ? mux_stage_4[174] : mux_stage_4[166];
	assign mux_stage_3[167] = (sel_3_reg0 == 1'b1) ? mux_stage_4[175] : mux_stage_4[167];
	assign mux_stage_3[168] = (sel_3_reg0 == 1'b1) ? mux_stage_4[176] : mux_stage_4[168];
	assign mux_stage_3[169] = (sel_3_reg0 == 1'b1) ? mux_stage_4[177] : mux_stage_4[169];
	assign mux_stage_3[170] = (sel_3_reg0 == 1'b1) ? mux_stage_4[178] : mux_stage_4[170];
	assign mux_stage_3[171] = (sel_3_reg0 == 1'b1) ? mux_stage_4[179] : mux_stage_4[171];
	assign mux_stage_3[172] = (sel_3_reg0 == 1'b1) ? mux_stage_4[180] : mux_stage_4[172];
	assign mux_stage_3[173] = (sel_3_reg0 == 1'b1) ? mux_stage_4[181] : mux_stage_4[173];
	assign mux_stage_3[174] = (sel_3_reg0 == 1'b1) ? mux_stage_4[182] : mux_stage_4[174];
	assign mux_stage_3[175] = (sel_3_reg0 == 1'b1) ? mux_stage_4[183] : mux_stage_4[175];
	assign mux_stage_3[176] = (sel_3_reg0 == 1'b1) ? mux_stage_4[184] : mux_stage_4[176];
	assign mux_stage_3[177] = (sel_3_reg0 == 1'b1) ? mux_stage_4[185] : mux_stage_4[177];
	assign mux_stage_3[178] = (sel_3_reg0 == 1'b1) ? mux_stage_4[186] : mux_stage_4[178];
	assign mux_stage_3[179] = (sel_3_reg0 == 1'b1) ? mux_stage_4[187] : mux_stage_4[179];
	assign mux_stage_3[180] = (sel_3_reg0 == 1'b1) ? mux_stage_4[188] : mux_stage_4[180];
	assign mux_stage_3[181] = (sel_3_reg0 == 1'b1) ? mux_stage_4[189] : mux_stage_4[181];
	assign mux_stage_3[182] = (sel_3_reg0 == 1'b1) ? mux_stage_4[190] : mux_stage_4[182];
	assign mux_stage_3[183] = (sel_3_reg0 == 1'b1) ? mux_stage_4[191] : mux_stage_4[183];
	assign mux_stage_3[184] = (sel_3_reg0 == 1'b1) ? mux_stage_4[192] : mux_stage_4[184];
	assign mux_stage_3[185] = (sel_3_reg0 == 1'b1) ? mux_stage_4[193] : mux_stage_4[185];
	assign mux_stage_3[186] = (sel_3_reg0 == 1'b1) ? mux_stage_4[194] : mux_stage_4[186];
	assign mux_stage_3[187] = (sel_3_reg0 == 1'b1) ? mux_stage_4[195] : mux_stage_4[187];
	assign mux_stage_3[188] = (sel_3_reg0 == 1'b1) ? mux_stage_4[196] : mux_stage_4[188];
	assign mux_stage_3[189] = (sel_3_reg0 == 1'b1) ? mux_stage_4[197] : mux_stage_4[189];
	assign mux_stage_3[190] = (sel_3_reg0 == 1'b1) ? mux_stage_4[198] : mux_stage_4[190];
	assign mux_stage_3[191] = (sel_3_reg0 == 1'b1) ? mux_stage_4[199] : mux_stage_4[191];
	assign mux_stage_3[192] = (sel_3_reg0 == 1'b1) ? mux_stage_4[200] : mux_stage_4[192];
	assign mux_stage_3[193] = (sel_3_reg0 == 1'b1) ? mux_stage_4[201] : mux_stage_4[193];
	assign mux_stage_3[194] = (sel_3_reg0 == 1'b1) ? mux_stage_4[202] : mux_stage_4[194];
	assign mux_stage_3[195] = (sel_3_reg0 == 1'b1) ? mux_stage_4[203] : mux_stage_4[195];
	assign mux_stage_3[196] = (sel_3_reg0 == 1'b1) ? mux_stage_4[204] : mux_stage_4[196];
	assign mux_stage_3[197] = (sel_3_reg0 == 1'b1) ? mux_stage_4[205] : mux_stage_4[197];
	assign mux_stage_3[198] = (sel_3_reg0 == 1'b1) ? mux_stage_4[206] : mux_stage_4[198];
	assign mux_stage_3[199] = (sel_3_reg0 == 1'b1) ? mux_stage_4[207] : mux_stage_4[199];
	assign mux_stage_3[200] = (sel_3_reg0 == 1'b1) ? mux_stage_4[208] : mux_stage_4[200];
	assign mux_stage_3[201] = (sel_3_reg0 == 1'b1) ? mux_stage_4[209] : mux_stage_4[201];
	assign mux_stage_3[202] = (sel_3_reg0 == 1'b1) ? mux_stage_4[210] : mux_stage_4[202];
	assign mux_stage_3[203] = (sel_3_reg0 == 1'b1) ? mux_stage_4[211] : mux_stage_4[203];
	assign mux_stage_3[204] = (sel_3_reg0 == 1'b1) ? mux_stage_4[212] : mux_stage_4[204];
	assign mux_stage_3[205] = (sel_3_reg0 == 1'b1) ? mux_stage_4[213] : mux_stage_4[205];
	assign mux_stage_3[206] = (sel_3_reg0 == 1'b1) ? mux_stage_4[214] : mux_stage_4[206];
	assign mux_stage_3[207] = (sel_3_reg0 == 1'b1) ? mux_stage_4[215] : mux_stage_4[207];
	assign mux_stage_3[208] = (sel_3_reg0 == 1'b1) ? mux_stage_4[216] : mux_stage_4[208];
	assign mux_stage_3[209] = (sel_3_reg0 == 1'b1) ? mux_stage_4[217] : mux_stage_4[209];
	assign mux_stage_3[210] = (sel_3_reg0 == 1'b1) ? mux_stage_4[218] : mux_stage_4[210];
	assign mux_stage_3[211] = (sel_3_reg0 == 1'b1) ? mux_stage_4[219] : mux_stage_4[211];
	assign mux_stage_3[212] = (sel_3_reg0 == 1'b1) ? mux_stage_4[220] : mux_stage_4[212];
	assign mux_stage_3[213] = (sel_3_reg0 == 1'b1) ? mux_stage_4[221] : mux_stage_4[213];
	assign mux_stage_3[214] = (sel_3_reg0 == 1'b1) ? mux_stage_4[222] : mux_stage_4[214];
	assign mux_stage_3[215] = (sel_3_reg0 == 1'b1) ? mux_stage_4[223] : mux_stage_4[215];
	assign mux_stage_3[216] = (sel_3_reg0 == 1'b1) ? mux_stage_4[224] : mux_stage_4[216];
	assign mux_stage_3[217] = (sel_3_reg0 == 1'b1) ? mux_stage_4[225] : mux_stage_4[217];
	assign mux_stage_3[218] = (sel_3_reg0 == 1'b1) ? mux_stage_4[226] : mux_stage_4[218];
	assign mux_stage_3[219] = (sel_3_reg0 == 1'b1) ? mux_stage_4[227] : mux_stage_4[219];
	assign mux_stage_3[220] = (sel_3_reg0 == 1'b1) ? mux_stage_4[228] : mux_stage_4[220];
	assign mux_stage_3[221] = (sel_3_reg0 == 1'b1) ? mux_stage_4[229] : mux_stage_4[221];
	assign mux_stage_3[222] = (sel_3_reg0 == 1'b1) ? mux_stage_4[230] : mux_stage_4[222];
	assign mux_stage_3[223] = (sel_3_reg0 == 1'b1) ? mux_stage_4[231] : mux_stage_4[223];
	assign mux_stage_3[224] = (sel_3_reg0 == 1'b1) ? mux_stage_4[232] : mux_stage_4[224];
	assign mux_stage_3[225] = (sel_3_reg0 == 1'b1) ? mux_stage_4[233] : mux_stage_4[225];
	assign mux_stage_3[226] = (sel_3_reg0 == 1'b1) ? mux_stage_4[234] : mux_stage_4[226];
	assign mux_stage_3[227] = (sel_3_reg0 == 1'b1) ? mux_stage_4[235] : mux_stage_4[227];
	assign mux_stage_3[228] = (sel_3_reg0 == 1'b1) ? mux_stage_4[236] : mux_stage_4[228];
	assign mux_stage_3[229] = (sel_3_reg0 == 1'b1) ? mux_stage_4[237] : mux_stage_4[229];
	assign mux_stage_3[230] = (sel_3_reg0 == 1'b1) ? mux_stage_4[238] : mux_stage_4[230];
	assign mux_stage_3[231] = (sel_3_reg0 == 1'b1) ? sw_in_239_reg0 : mux_stage_4[231];
	assign mux_stage_3[232] = (sel_3_reg0 == 1'b1) ? sw_in_240_reg0 : mux_stage_4[232];
	assign mux_stage_3[233] = (sel_3_reg0 == 1'b1) ? sw_in_241_reg0 : mux_stage_4[233];
	assign mux_stage_3[234] = (sel_3_reg0 == 1'b1) ? sw_in_242_reg0 : mux_stage_4[234];
	assign mux_stage_3[235] = (sel_3_reg0 == 1'b1) ? sw_in_243_reg0 : mux_stage_4[235];
	assign mux_stage_3[236] = (sel_3_reg0 == 1'b1) ? sw_in_244_reg0 : mux_stage_4[236];
	assign mux_stage_3[237] = (sel_3_reg0 == 1'b1) ? sw_in_245_reg0 : mux_stage_4[237];
	assign mux_stage_3[238] = (sel_3_reg0 == 1'b1) ? sw_in_246_reg0 : mux_stage_4[238];
	assign mux_stage_3[239] = (sel_3_reg0 == 1'b1) ? sw_in_247_reg0 : sw_in_239_reg0;
	assign mux_stage_3[240] = (sel_3_reg0 == 1'b1) ? sw_in_248_reg0 : sw_in_240_reg0;
	assign mux_stage_3[241] = (sel_3_reg0 == 1'b1) ? sw_in_249_reg0 : sw_in_241_reg0;
	assign mux_stage_3[242] = (sel_3_reg0 == 1'b1) ? sw_in_250_reg0 : sw_in_242_reg0;
	assign mux_stage_3[243] = (sel_3_reg0 == 1'b1) ? sw_in_251_reg0 : sw_in_243_reg0;
	assign mux_stage_3[244] = (sel_3_reg0 == 1'b1) ? sw_in_252_reg0 : sw_in_244_reg0;
	assign mux_stage_3[245] = (sel_3_reg0 == 1'b1) ? sw_in_253_reg0 : sw_in_245_reg0;
	assign mux_stage_3[246] = (sel_3_reg0 == 1'b1) ? sw_in_254_reg0 : sw_in_246_reg0;


	reg sel_2_reg0;
	always @(posedge sys_clk) begin if(!rstn) sel_2_reg0 <= 0; else sel_2_reg0 <= sel[2]; end	

	// Multiplexer Stage 2
	wire [250:0] mux_stage_2;
	assign mux_stage_2[0] = (sel_2_reg0 == 1'b1) ? mux_stage_3[4] : mux_stage_3[0];
	assign mux_stage_2[1] = (sel_2_reg0 == 1'b1) ? mux_stage_3[5] : mux_stage_3[1];
	assign mux_stage_2[2] = (sel_2_reg0 == 1'b1) ? mux_stage_3[6] : mux_stage_3[2];
	assign mux_stage_2[3] = (sel_2_reg0 == 1'b1) ? mux_stage_3[7] : mux_stage_3[3];
	assign mux_stage_2[4] = (sel_2_reg0 == 1'b1) ? mux_stage_3[8] : mux_stage_3[4];
	assign mux_stage_2[5] = (sel_2_reg0 == 1'b1) ? mux_stage_3[9] : mux_stage_3[5];
	assign mux_stage_2[6] = (sel_2_reg0 == 1'b1) ? mux_stage_3[10] : mux_stage_3[6];
	assign mux_stage_2[7] = (sel_2_reg0 == 1'b1) ? mux_stage_3[11] : mux_stage_3[7];
	assign mux_stage_2[8] = (sel_2_reg0 == 1'b1) ? mux_stage_3[12] : mux_stage_3[8];
	assign mux_stage_2[9] = (sel_2_reg0 == 1'b1) ? mux_stage_3[13] : mux_stage_3[9];
	assign mux_stage_2[10] = (sel_2_reg0 == 1'b1) ? mux_stage_3[14] : mux_stage_3[10];
	assign mux_stage_2[11] = (sel_2_reg0 == 1'b1) ? mux_stage_3[15] : mux_stage_3[11];
	assign mux_stage_2[12] = (sel_2_reg0 == 1'b1) ? mux_stage_3[16] : mux_stage_3[12];
	assign mux_stage_2[13] = (sel_2_reg0 == 1'b1) ? mux_stage_3[17] : mux_stage_3[13];
	assign mux_stage_2[14] = (sel_2_reg0 == 1'b1) ? mux_stage_3[18] : mux_stage_3[14];
	assign mux_stage_2[15] = (sel_2_reg0 == 1'b1) ? mux_stage_3[19] : mux_stage_3[15];
	assign mux_stage_2[16] = (sel_2_reg0 == 1'b1) ? mux_stage_3[20] : mux_stage_3[16];
	assign mux_stage_2[17] = (sel_2_reg0 == 1'b1) ? mux_stage_3[21] : mux_stage_3[17];
	assign mux_stage_2[18] = (sel_2_reg0 == 1'b1) ? mux_stage_3[22] : mux_stage_3[18];
	assign mux_stage_2[19] = (sel_2_reg0 == 1'b1) ? mux_stage_3[23] : mux_stage_3[19];
	assign mux_stage_2[20] = (sel_2_reg0 == 1'b1) ? mux_stage_3[24] : mux_stage_3[20];
	assign mux_stage_2[21] = (sel_2_reg0 == 1'b1) ? mux_stage_3[25] : mux_stage_3[21];
	assign mux_stage_2[22] = (sel_2_reg0 == 1'b1) ? mux_stage_3[26] : mux_stage_3[22];
	assign mux_stage_2[23] = (sel_2_reg0 == 1'b1) ? mux_stage_3[27] : mux_stage_3[23];
	assign mux_stage_2[24] = (sel_2_reg0 == 1'b1) ? mux_stage_3[28] : mux_stage_3[24];
	assign mux_stage_2[25] = (sel_2_reg0 == 1'b1) ? mux_stage_3[29] : mux_stage_3[25];
	assign mux_stage_2[26] = (sel_2_reg0 == 1'b1) ? mux_stage_3[30] : mux_stage_3[26];
	assign mux_stage_2[27] = (sel_2_reg0 == 1'b1) ? mux_stage_3[31] : mux_stage_3[27];
	assign mux_stage_2[28] = (sel_2_reg0 == 1'b1) ? mux_stage_3[32] : mux_stage_3[28];
	assign mux_stage_2[29] = (sel_2_reg0 == 1'b1) ? mux_stage_3[33] : mux_stage_3[29];
	assign mux_stage_2[30] = (sel_2_reg0 == 1'b1) ? mux_stage_3[34] : mux_stage_3[30];
	assign mux_stage_2[31] = (sel_2_reg0 == 1'b1) ? mux_stage_3[35] : mux_stage_3[31];
	assign mux_stage_2[32] = (sel_2_reg0 == 1'b1) ? mux_stage_3[36] : mux_stage_3[32];
	assign mux_stage_2[33] = (sel_2_reg0 == 1'b1) ? mux_stage_3[37] : mux_stage_3[33];
	assign mux_stage_2[34] = (sel_2_reg0 == 1'b1) ? mux_stage_3[38] : mux_stage_3[34];
	assign mux_stage_2[35] = (sel_2_reg0 == 1'b1) ? mux_stage_3[39] : mux_stage_3[35];
	assign mux_stage_2[36] = (sel_2_reg0 == 1'b1) ? mux_stage_3[40] : mux_stage_3[36];
	assign mux_stage_2[37] = (sel_2_reg0 == 1'b1) ? mux_stage_3[41] : mux_stage_3[37];
	assign mux_stage_2[38] = (sel_2_reg0 == 1'b1) ? mux_stage_3[42] : mux_stage_3[38];
	assign mux_stage_2[39] = (sel_2_reg0 == 1'b1) ? mux_stage_3[43] : mux_stage_3[39];
	assign mux_stage_2[40] = (sel_2_reg0 == 1'b1) ? mux_stage_3[44] : mux_stage_3[40];
	assign mux_stage_2[41] = (sel_2_reg0 == 1'b1) ? mux_stage_3[45] : mux_stage_3[41];
	assign mux_stage_2[42] = (sel_2_reg0 == 1'b1) ? mux_stage_3[46] : mux_stage_3[42];
	assign mux_stage_2[43] = (sel_2_reg0 == 1'b1) ? mux_stage_3[47] : mux_stage_3[43];
	assign mux_stage_2[44] = (sel_2_reg0 == 1'b1) ? mux_stage_3[48] : mux_stage_3[44];
	assign mux_stage_2[45] = (sel_2_reg0 == 1'b1) ? mux_stage_3[49] : mux_stage_3[45];
	assign mux_stage_2[46] = (sel_2_reg0 == 1'b1) ? mux_stage_3[50] : mux_stage_3[46];
	assign mux_stage_2[47] = (sel_2_reg0 == 1'b1) ? mux_stage_3[51] : mux_stage_3[47];
	assign mux_stage_2[48] = (sel_2_reg0 == 1'b1) ? mux_stage_3[52] : mux_stage_3[48];
	assign mux_stage_2[49] = (sel_2_reg0 == 1'b1) ? mux_stage_3[53] : mux_stage_3[49];
	assign mux_stage_2[50] = (sel_2_reg0 == 1'b1) ? mux_stage_3[54] : mux_stage_3[50];
	assign mux_stage_2[51] = (sel_2_reg0 == 1'b1) ? mux_stage_3[55] : mux_stage_3[51];
	assign mux_stage_2[52] = (sel_2_reg0 == 1'b1) ? mux_stage_3[56] : mux_stage_3[52];
	assign mux_stage_2[53] = (sel_2_reg0 == 1'b1) ? mux_stage_3[57] : mux_stage_3[53];
	assign mux_stage_2[54] = (sel_2_reg0 == 1'b1) ? mux_stage_3[58] : mux_stage_3[54];
	assign mux_stage_2[55] = (sel_2_reg0 == 1'b1) ? mux_stage_3[59] : mux_stage_3[55];
	assign mux_stage_2[56] = (sel_2_reg0 == 1'b1) ? mux_stage_3[60] : mux_stage_3[56];
	assign mux_stage_2[57] = (sel_2_reg0 == 1'b1) ? mux_stage_3[61] : mux_stage_3[57];
	assign mux_stage_2[58] = (sel_2_reg0 == 1'b1) ? mux_stage_3[62] : mux_stage_3[58];
	assign mux_stage_2[59] = (sel_2_reg0 == 1'b1) ? mux_stage_3[63] : mux_stage_3[59];
	assign mux_stage_2[60] = (sel_2_reg0 == 1'b1) ? mux_stage_3[64] : mux_stage_3[60];
	assign mux_stage_2[61] = (sel_2_reg0 == 1'b1) ? mux_stage_3[65] : mux_stage_3[61];
	assign mux_stage_2[62] = (sel_2_reg0 == 1'b1) ? mux_stage_3[66] : mux_stage_3[62];
	assign mux_stage_2[63] = (sel_2_reg0 == 1'b1) ? mux_stage_3[67] : mux_stage_3[63];
	assign mux_stage_2[64] = (sel_2_reg0 == 1'b1) ? mux_stage_3[68] : mux_stage_3[64];
	assign mux_stage_2[65] = (sel_2_reg0 == 1'b1) ? mux_stage_3[69] : mux_stage_3[65];
	assign mux_stage_2[66] = (sel_2_reg0 == 1'b1) ? mux_stage_3[70] : mux_stage_3[66];
	assign mux_stage_2[67] = (sel_2_reg0 == 1'b1) ? mux_stage_3[71] : mux_stage_3[67];
	assign mux_stage_2[68] = (sel_2_reg0 == 1'b1) ? mux_stage_3[72] : mux_stage_3[68];
	assign mux_stage_2[69] = (sel_2_reg0 == 1'b1) ? mux_stage_3[73] : mux_stage_3[69];
	assign mux_stage_2[70] = (sel_2_reg0 == 1'b1) ? mux_stage_3[74] : mux_stage_3[70];
	assign mux_stage_2[71] = (sel_2_reg0 == 1'b1) ? mux_stage_3[75] : mux_stage_3[71];
	assign mux_stage_2[72] = (sel_2_reg0 == 1'b1) ? mux_stage_3[76] : mux_stage_3[72];
	assign mux_stage_2[73] = (sel_2_reg0 == 1'b1) ? mux_stage_3[77] : mux_stage_3[73];
	assign mux_stage_2[74] = (sel_2_reg0 == 1'b1) ? mux_stage_3[78] : mux_stage_3[74];
	assign mux_stage_2[75] = (sel_2_reg0 == 1'b1) ? mux_stage_3[79] : mux_stage_3[75];
	assign mux_stage_2[76] = (sel_2_reg0 == 1'b1) ? mux_stage_3[80] : mux_stage_3[76];
	assign mux_stage_2[77] = (sel_2_reg0 == 1'b1) ? mux_stage_3[81] : mux_stage_3[77];
	assign mux_stage_2[78] = (sel_2_reg0 == 1'b1) ? mux_stage_3[82] : mux_stage_3[78];
	assign mux_stage_2[79] = (sel_2_reg0 == 1'b1) ? mux_stage_3[83] : mux_stage_3[79];
	assign mux_stage_2[80] = (sel_2_reg0 == 1'b1) ? mux_stage_3[84] : mux_stage_3[80];
	assign mux_stage_2[81] = (sel_2_reg0 == 1'b1) ? mux_stage_3[85] : mux_stage_3[81];
	assign mux_stage_2[82] = (sel_2_reg0 == 1'b1) ? mux_stage_3[86] : mux_stage_3[82];
	assign mux_stage_2[83] = (sel_2_reg0 == 1'b1) ? mux_stage_3[87] : mux_stage_3[83];
	assign mux_stage_2[84] = (sel_2_reg0 == 1'b1) ? mux_stage_3[88] : mux_stage_3[84];
	assign mux_stage_2[85] = (sel_2_reg0 == 1'b1) ? mux_stage_3[89] : mux_stage_3[85];
	assign mux_stage_2[86] = (sel_2_reg0 == 1'b1) ? mux_stage_3[90] : mux_stage_3[86];
	assign mux_stage_2[87] = (sel_2_reg0 == 1'b1) ? mux_stage_3[91] : mux_stage_3[87];
	assign mux_stage_2[88] = (sel_2_reg0 == 1'b1) ? mux_stage_3[92] : mux_stage_3[88];
	assign mux_stage_2[89] = (sel_2_reg0 == 1'b1) ? mux_stage_3[93] : mux_stage_3[89];
	assign mux_stage_2[90] = (sel_2_reg0 == 1'b1) ? mux_stage_3[94] : mux_stage_3[90];
	assign mux_stage_2[91] = (sel_2_reg0 == 1'b1) ? mux_stage_3[95] : mux_stage_3[91];
	assign mux_stage_2[92] = (sel_2_reg0 == 1'b1) ? mux_stage_3[96] : mux_stage_3[92];
	assign mux_stage_2[93] = (sel_2_reg0 == 1'b1) ? mux_stage_3[97] : mux_stage_3[93];
	assign mux_stage_2[94] = (sel_2_reg0 == 1'b1) ? mux_stage_3[98] : mux_stage_3[94];
	assign mux_stage_2[95] = (sel_2_reg0 == 1'b1) ? mux_stage_3[99] : mux_stage_3[95];
	assign mux_stage_2[96] = (sel_2_reg0 == 1'b1) ? mux_stage_3[100] : mux_stage_3[96];
	assign mux_stage_2[97] = (sel_2_reg0 == 1'b1) ? mux_stage_3[101] : mux_stage_3[97];
	assign mux_stage_2[98] = (sel_2_reg0 == 1'b1) ? mux_stage_3[102] : mux_stage_3[98];
	assign mux_stage_2[99] = (sel_2_reg0 == 1'b1) ? mux_stage_3[103] : mux_stage_3[99];
	assign mux_stage_2[100] = (sel_2_reg0 == 1'b1) ? mux_stage_3[104] : mux_stage_3[100];
	assign mux_stage_2[101] = (sel_2_reg0 == 1'b1) ? mux_stage_3[105] : mux_stage_3[101];
	assign mux_stage_2[102] = (sel_2_reg0 == 1'b1) ? mux_stage_3[106] : mux_stage_3[102];
	assign mux_stage_2[103] = (sel_2_reg0 == 1'b1) ? mux_stage_3[107] : mux_stage_3[103];
	assign mux_stage_2[104] = (sel_2_reg0 == 1'b1) ? mux_stage_3[108] : mux_stage_3[104];
	assign mux_stage_2[105] = (sel_2_reg0 == 1'b1) ? mux_stage_3[109] : mux_stage_3[105];
	assign mux_stage_2[106] = (sel_2_reg0 == 1'b1) ? mux_stage_3[110] : mux_stage_3[106];
	assign mux_stage_2[107] = (sel_2_reg0 == 1'b1) ? mux_stage_3[111] : mux_stage_3[107];
	assign mux_stage_2[108] = (sel_2_reg0 == 1'b1) ? mux_stage_3[112] : mux_stage_3[108];
	assign mux_stage_2[109] = (sel_2_reg0 == 1'b1) ? mux_stage_3[113] : mux_stage_3[109];
	assign mux_stage_2[110] = (sel_2_reg0 == 1'b1) ? mux_stage_3[114] : mux_stage_3[110];
	assign mux_stage_2[111] = (sel_2_reg0 == 1'b1) ? mux_stage_3[115] : mux_stage_3[111];
	assign mux_stage_2[112] = (sel_2_reg0 == 1'b1) ? mux_stage_3[116] : mux_stage_3[112];
	assign mux_stage_2[113] = (sel_2_reg0 == 1'b1) ? mux_stage_3[117] : mux_stage_3[113];
	assign mux_stage_2[114] = (sel_2_reg0 == 1'b1) ? mux_stage_3[118] : mux_stage_3[114];
	assign mux_stage_2[115] = (sel_2_reg0 == 1'b1) ? mux_stage_3[119] : mux_stage_3[115];
	assign mux_stage_2[116] = (sel_2_reg0 == 1'b1) ? mux_stage_3[120] : mux_stage_3[116];
	assign mux_stage_2[117] = (sel_2_reg0 == 1'b1) ? mux_stage_3[121] : mux_stage_3[117];
	assign mux_stage_2[118] = (sel_2_reg0 == 1'b1) ? mux_stage_3[122] : mux_stage_3[118];
	assign mux_stage_2[119] = (sel_2_reg0 == 1'b1) ? mux_stage_3[123] : mux_stage_3[119];
	assign mux_stage_2[120] = (sel_2_reg0 == 1'b1) ? mux_stage_3[124] : mux_stage_3[120];
	assign mux_stage_2[121] = (sel_2_reg0 == 1'b1) ? mux_stage_3[125] : mux_stage_3[121];
	assign mux_stage_2[122] = (sel_2_reg0 == 1'b1) ? mux_stage_3[126] : mux_stage_3[122];
	assign mux_stage_2[123] = (sel_2_reg0 == 1'b1) ? mux_stage_3[127] : mux_stage_3[123];
	assign mux_stage_2[124] = (sel_2_reg0 == 1'b1) ? mux_stage_3[128] : mux_stage_3[124];
	assign mux_stage_2[125] = (sel_2_reg0 == 1'b1) ? mux_stage_3[129] : mux_stage_3[125];
	assign mux_stage_2[126] = (sel_2_reg0 == 1'b1) ? mux_stage_3[130] : mux_stage_3[126];
	assign mux_stage_2[127] = (sel_2_reg0 == 1'b1) ? mux_stage_3[131] : mux_stage_3[127];
	assign mux_stage_2[128] = (sel_2_reg0 == 1'b1) ? mux_stage_3[132] : mux_stage_3[128];
	assign mux_stage_2[129] = (sel_2_reg0 == 1'b1) ? mux_stage_3[133] : mux_stage_3[129];
	assign mux_stage_2[130] = (sel_2_reg0 == 1'b1) ? mux_stage_3[134] : mux_stage_3[130];
	assign mux_stage_2[131] = (sel_2_reg0 == 1'b1) ? mux_stage_3[135] : mux_stage_3[131];
	assign mux_stage_2[132] = (sel_2_reg0 == 1'b1) ? mux_stage_3[136] : mux_stage_3[132];
	assign mux_stage_2[133] = (sel_2_reg0 == 1'b1) ? mux_stage_3[137] : mux_stage_3[133];
	assign mux_stage_2[134] = (sel_2_reg0 == 1'b1) ? mux_stage_3[138] : mux_stage_3[134];
	assign mux_stage_2[135] = (sel_2_reg0 == 1'b1) ? mux_stage_3[139] : mux_stage_3[135];
	assign mux_stage_2[136] = (sel_2_reg0 == 1'b1) ? mux_stage_3[140] : mux_stage_3[136];
	assign mux_stage_2[137] = (sel_2_reg0 == 1'b1) ? mux_stage_3[141] : mux_stage_3[137];
	assign mux_stage_2[138] = (sel_2_reg0 == 1'b1) ? mux_stage_3[142] : mux_stage_3[138];
	assign mux_stage_2[139] = (sel_2_reg0 == 1'b1) ? mux_stage_3[143] : mux_stage_3[139];
	assign mux_stage_2[140] = (sel_2_reg0 == 1'b1) ? mux_stage_3[144] : mux_stage_3[140];
	assign mux_stage_2[141] = (sel_2_reg0 == 1'b1) ? mux_stage_3[145] : mux_stage_3[141];
	assign mux_stage_2[142] = (sel_2_reg0 == 1'b1) ? mux_stage_3[146] : mux_stage_3[142];
	assign mux_stage_2[143] = (sel_2_reg0 == 1'b1) ? mux_stage_3[147] : mux_stage_3[143];
	assign mux_stage_2[144] = (sel_2_reg0 == 1'b1) ? mux_stage_3[148] : mux_stage_3[144];
	assign mux_stage_2[145] = (sel_2_reg0 == 1'b1) ? mux_stage_3[149] : mux_stage_3[145];
	assign mux_stage_2[146] = (sel_2_reg0 == 1'b1) ? mux_stage_3[150] : mux_stage_3[146];
	assign mux_stage_2[147] = (sel_2_reg0 == 1'b1) ? mux_stage_3[151] : mux_stage_3[147];
	assign mux_stage_2[148] = (sel_2_reg0 == 1'b1) ? mux_stage_3[152] : mux_stage_3[148];
	assign mux_stage_2[149] = (sel_2_reg0 == 1'b1) ? mux_stage_3[153] : mux_stage_3[149];
	assign mux_stage_2[150] = (sel_2_reg0 == 1'b1) ? mux_stage_3[154] : mux_stage_3[150];
	assign mux_stage_2[151] = (sel_2_reg0 == 1'b1) ? mux_stage_3[155] : mux_stage_3[151];
	assign mux_stage_2[152] = (sel_2_reg0 == 1'b1) ? mux_stage_3[156] : mux_stage_3[152];
	assign mux_stage_2[153] = (sel_2_reg0 == 1'b1) ? mux_stage_3[157] : mux_stage_3[153];
	assign mux_stage_2[154] = (sel_2_reg0 == 1'b1) ? mux_stage_3[158] : mux_stage_3[154];
	assign mux_stage_2[155] = (sel_2_reg0 == 1'b1) ? mux_stage_3[159] : mux_stage_3[155];
	assign mux_stage_2[156] = (sel_2_reg0 == 1'b1) ? mux_stage_3[160] : mux_stage_3[156];
	assign mux_stage_2[157] = (sel_2_reg0 == 1'b1) ? mux_stage_3[161] : mux_stage_3[157];
	assign mux_stage_2[158] = (sel_2_reg0 == 1'b1) ? mux_stage_3[162] : mux_stage_3[158];
	assign mux_stage_2[159] = (sel_2_reg0 == 1'b1) ? mux_stage_3[163] : mux_stage_3[159];
	assign mux_stage_2[160] = (sel_2_reg0 == 1'b1) ? mux_stage_3[164] : mux_stage_3[160];
	assign mux_stage_2[161] = (sel_2_reg0 == 1'b1) ? mux_stage_3[165] : mux_stage_3[161];
	assign mux_stage_2[162] = (sel_2_reg0 == 1'b1) ? mux_stage_3[166] : mux_stage_3[162];
	assign mux_stage_2[163] = (sel_2_reg0 == 1'b1) ? mux_stage_3[167] : mux_stage_3[163];
	assign mux_stage_2[164] = (sel_2_reg0 == 1'b1) ? mux_stage_3[168] : mux_stage_3[164];
	assign mux_stage_2[165] = (sel_2_reg0 == 1'b1) ? mux_stage_3[169] : mux_stage_3[165];
	assign mux_stage_2[166] = (sel_2_reg0 == 1'b1) ? mux_stage_3[170] : mux_stage_3[166];
	assign mux_stage_2[167] = (sel_2_reg0 == 1'b1) ? mux_stage_3[171] : mux_stage_3[167];
	assign mux_stage_2[168] = (sel_2_reg0 == 1'b1) ? mux_stage_3[172] : mux_stage_3[168];
	assign mux_stage_2[169] = (sel_2_reg0 == 1'b1) ? mux_stage_3[173] : mux_stage_3[169];
	assign mux_stage_2[170] = (sel_2_reg0 == 1'b1) ? mux_stage_3[174] : mux_stage_3[170];
	assign mux_stage_2[171] = (sel_2_reg0 == 1'b1) ? mux_stage_3[175] : mux_stage_3[171];
	assign mux_stage_2[172] = (sel_2_reg0 == 1'b1) ? mux_stage_3[176] : mux_stage_3[172];
	assign mux_stage_2[173] = (sel_2_reg0 == 1'b1) ? mux_stage_3[177] : mux_stage_3[173];
	assign mux_stage_2[174] = (sel_2_reg0 == 1'b1) ? mux_stage_3[178] : mux_stage_3[174];
	assign mux_stage_2[175] = (sel_2_reg0 == 1'b1) ? mux_stage_3[179] : mux_stage_3[175];
	assign mux_stage_2[176] = (sel_2_reg0 == 1'b1) ? mux_stage_3[180] : mux_stage_3[176];
	assign mux_stage_2[177] = (sel_2_reg0 == 1'b1) ? mux_stage_3[181] : mux_stage_3[177];
	assign mux_stage_2[178] = (sel_2_reg0 == 1'b1) ? mux_stage_3[182] : mux_stage_3[178];
	assign mux_stage_2[179] = (sel_2_reg0 == 1'b1) ? mux_stage_3[183] : mux_stage_3[179];
	assign mux_stage_2[180] = (sel_2_reg0 == 1'b1) ? mux_stage_3[184] : mux_stage_3[180];
	assign mux_stage_2[181] = (sel_2_reg0 == 1'b1) ? mux_stage_3[185] : mux_stage_3[181];
	assign mux_stage_2[182] = (sel_2_reg0 == 1'b1) ? mux_stage_3[186] : mux_stage_3[182];
	assign mux_stage_2[183] = (sel_2_reg0 == 1'b1) ? mux_stage_3[187] : mux_stage_3[183];
	assign mux_stage_2[184] = (sel_2_reg0 == 1'b1) ? mux_stage_3[188] : mux_stage_3[184];
	assign mux_stage_2[185] = (sel_2_reg0 == 1'b1) ? mux_stage_3[189] : mux_stage_3[185];
	assign mux_stage_2[186] = (sel_2_reg0 == 1'b1) ? mux_stage_3[190] : mux_stage_3[186];
	assign mux_stage_2[187] = (sel_2_reg0 == 1'b1) ? mux_stage_3[191] : mux_stage_3[187];
	assign mux_stage_2[188] = (sel_2_reg0 == 1'b1) ? mux_stage_3[192] : mux_stage_3[188];
	assign mux_stage_2[189] = (sel_2_reg0 == 1'b1) ? mux_stage_3[193] : mux_stage_3[189];
	assign mux_stage_2[190] = (sel_2_reg0 == 1'b1) ? mux_stage_3[194] : mux_stage_3[190];
	assign mux_stage_2[191] = (sel_2_reg0 == 1'b1) ? mux_stage_3[195] : mux_stage_3[191];
	assign mux_stage_2[192] = (sel_2_reg0 == 1'b1) ? mux_stage_3[196] : mux_stage_3[192];
	assign mux_stage_2[193] = (sel_2_reg0 == 1'b1) ? mux_stage_3[197] : mux_stage_3[193];
	assign mux_stage_2[194] = (sel_2_reg0 == 1'b1) ? mux_stage_3[198] : mux_stage_3[194];
	assign mux_stage_2[195] = (sel_2_reg0 == 1'b1) ? mux_stage_3[199] : mux_stage_3[195];
	assign mux_stage_2[196] = (sel_2_reg0 == 1'b1) ? mux_stage_3[200] : mux_stage_3[196];
	assign mux_stage_2[197] = (sel_2_reg0 == 1'b1) ? mux_stage_3[201] : mux_stage_3[197];
	assign mux_stage_2[198] = (sel_2_reg0 == 1'b1) ? mux_stage_3[202] : mux_stage_3[198];
	assign mux_stage_2[199] = (sel_2_reg0 == 1'b1) ? mux_stage_3[203] : mux_stage_3[199];
	assign mux_stage_2[200] = (sel_2_reg0 == 1'b1) ? mux_stage_3[204] : mux_stage_3[200];
	assign mux_stage_2[201] = (sel_2_reg0 == 1'b1) ? mux_stage_3[205] : mux_stage_3[201];
	assign mux_stage_2[202] = (sel_2_reg0 == 1'b1) ? mux_stage_3[206] : mux_stage_3[202];
	assign mux_stage_2[203] = (sel_2_reg0 == 1'b1) ? mux_stage_3[207] : mux_stage_3[203];
	assign mux_stage_2[204] = (sel_2_reg0 == 1'b1) ? mux_stage_3[208] : mux_stage_3[204];
	assign mux_stage_2[205] = (sel_2_reg0 == 1'b1) ? mux_stage_3[209] : mux_stage_3[205];
	assign mux_stage_2[206] = (sel_2_reg0 == 1'b1) ? mux_stage_3[210] : mux_stage_3[206];
	assign mux_stage_2[207] = (sel_2_reg0 == 1'b1) ? mux_stage_3[211] : mux_stage_3[207];
	assign mux_stage_2[208] = (sel_2_reg0 == 1'b1) ? mux_stage_3[212] : mux_stage_3[208];
	assign mux_stage_2[209] = (sel_2_reg0 == 1'b1) ? mux_stage_3[213] : mux_stage_3[209];
	assign mux_stage_2[210] = (sel_2_reg0 == 1'b1) ? mux_stage_3[214] : mux_stage_3[210];
	assign mux_stage_2[211] = (sel_2_reg0 == 1'b1) ? mux_stage_3[215] : mux_stage_3[211];
	assign mux_stage_2[212] = (sel_2_reg0 == 1'b1) ? mux_stage_3[216] : mux_stage_3[212];
	assign mux_stage_2[213] = (sel_2_reg0 == 1'b1) ? mux_stage_3[217] : mux_stage_3[213];
	assign mux_stage_2[214] = (sel_2_reg0 == 1'b1) ? mux_stage_3[218] : mux_stage_3[214];
	assign mux_stage_2[215] = (sel_2_reg0 == 1'b1) ? mux_stage_3[219] : mux_stage_3[215];
	assign mux_stage_2[216] = (sel_2_reg0 == 1'b1) ? mux_stage_3[220] : mux_stage_3[216];
	assign mux_stage_2[217] = (sel_2_reg0 == 1'b1) ? mux_stage_3[221] : mux_stage_3[217];
	assign mux_stage_2[218] = (sel_2_reg0 == 1'b1) ? mux_stage_3[222] : mux_stage_3[218];
	assign mux_stage_2[219] = (sel_2_reg0 == 1'b1) ? mux_stage_3[223] : mux_stage_3[219];
	assign mux_stage_2[220] = (sel_2_reg0 == 1'b1) ? mux_stage_3[224] : mux_stage_3[220];
	assign mux_stage_2[221] = (sel_2_reg0 == 1'b1) ? mux_stage_3[225] : mux_stage_3[221];
	assign mux_stage_2[222] = (sel_2_reg0 == 1'b1) ? mux_stage_3[226] : mux_stage_3[222];
	assign mux_stage_2[223] = (sel_2_reg0 == 1'b1) ? mux_stage_3[227] : mux_stage_3[223];
	assign mux_stage_2[224] = (sel_2_reg0 == 1'b1) ? mux_stage_3[228] : mux_stage_3[224];
	assign mux_stage_2[225] = (sel_2_reg0 == 1'b1) ? mux_stage_3[229] : mux_stage_3[225];
	assign mux_stage_2[226] = (sel_2_reg0 == 1'b1) ? mux_stage_3[230] : mux_stage_3[226];
	assign mux_stage_2[227] = (sel_2_reg0 == 1'b1) ? mux_stage_3[231] : mux_stage_3[227];
	assign mux_stage_2[228] = (sel_2_reg0 == 1'b1) ? mux_stage_3[232] : mux_stage_3[228];
	assign mux_stage_2[229] = (sel_2_reg0 == 1'b1) ? mux_stage_3[233] : mux_stage_3[229];
	assign mux_stage_2[230] = (sel_2_reg0 == 1'b1) ? mux_stage_3[234] : mux_stage_3[230];
	assign mux_stage_2[231] = (sel_2_reg0 == 1'b1) ? mux_stage_3[235] : mux_stage_3[231];
	assign mux_stage_2[232] = (sel_2_reg0 == 1'b1) ? mux_stage_3[236] : mux_stage_3[232];
	assign mux_stage_2[233] = (sel_2_reg0 == 1'b1) ? mux_stage_3[237] : mux_stage_3[233];
	assign mux_stage_2[234] = (sel_2_reg0 == 1'b1) ? mux_stage_3[238] : mux_stage_3[234];
	assign mux_stage_2[235] = (sel_2_reg0 == 1'b1) ? mux_stage_3[239] : mux_stage_3[235];
	assign mux_stage_2[236] = (sel_2_reg0 == 1'b1) ? mux_stage_3[240] : mux_stage_3[236];
	assign mux_stage_2[237] = (sel_2_reg0 == 1'b1) ? mux_stage_3[241] : mux_stage_3[237];
	assign mux_stage_2[238] = (sel_2_reg0 == 1'b1) ? mux_stage_3[242] : mux_stage_3[238];
	assign mux_stage_2[239] = (sel_2_reg0 == 1'b1) ? mux_stage_3[243] : mux_stage_3[239];
	assign mux_stage_2[240] = (sel_2_reg0 == 1'b1) ? mux_stage_3[244] : mux_stage_3[240];
	assign mux_stage_2[241] = (sel_2_reg0 == 1'b1) ? mux_stage_3[245] : mux_stage_3[241];
	assign mux_stage_2[242] = (sel_2_reg0 == 1'b1) ? mux_stage_3[246] : mux_stage_3[242];
	assign mux_stage_2[243] = (sel_2_reg0 == 1'b1) ? sw_in_247_reg0 : mux_stage_3[243];
	assign mux_stage_2[244] = (sel_2_reg0 == 1'b1) ? sw_in_248_reg0 : mux_stage_3[244];
	assign mux_stage_2[245] = (sel_2_reg0 == 1'b1) ? sw_in_249_reg0 : mux_stage_3[245];
	assign mux_stage_2[246] = (sel_2_reg0 == 1'b1) ? sw_in_250_reg0 : mux_stage_3[246];
	assign mux_stage_2[247] = (sel_2_reg0 == 1'b1) ? sw_in_251_reg0 : sw_in_247_reg0;
	assign mux_stage_2[248] = (sel_2_reg0 == 1'b1) ? sw_in_252_reg0 : sw_in_248_reg0;
	assign mux_stage_2[249] = (sel_2_reg0 == 1'b1) ? sw_in_253_reg0 : sw_in_249_reg0;
	assign mux_stage_2[250] = (sel_2_reg0 == 1'b1) ? sw_in_254_reg0 : sw_in_250_reg0;


	reg sel_1_reg0;
	always @(posedge sys_clk) begin if(!rstn) sel_1_reg0 <= 0; else sel_1_reg0 <= sel[1]; end	

	// Multiplexer Stage 1
	wire [252:0] mux_stage_1;
	assign mux_stage_1[0] = (sel_1_reg0 == 1'b1) ? mux_stage_2[2] : mux_stage_2[0];
	assign mux_stage_1[1] = (sel_1_reg0 == 1'b1) ? mux_stage_2[3] : mux_stage_2[1];
	assign mux_stage_1[2] = (sel_1_reg0 == 1'b1) ? mux_stage_2[4] : mux_stage_2[2];
	assign mux_stage_1[3] = (sel_1_reg0 == 1'b1) ? mux_stage_2[5] : mux_stage_2[3];
	assign mux_stage_1[4] = (sel_1_reg0 == 1'b1) ? mux_stage_2[6] : mux_stage_2[4];
	assign mux_stage_1[5] = (sel_1_reg0 == 1'b1) ? mux_stage_2[7] : mux_stage_2[5];
	assign mux_stage_1[6] = (sel_1_reg0 == 1'b1) ? mux_stage_2[8] : mux_stage_2[6];
	assign mux_stage_1[7] = (sel_1_reg0 == 1'b1) ? mux_stage_2[9] : mux_stage_2[7];
	assign mux_stage_1[8] = (sel_1_reg0 == 1'b1) ? mux_stage_2[10] : mux_stage_2[8];
	assign mux_stage_1[9] = (sel_1_reg0 == 1'b1) ? mux_stage_2[11] : mux_stage_2[9];
	assign mux_stage_1[10] = (sel_1_reg0 == 1'b1) ? mux_stage_2[12] : mux_stage_2[10];
	assign mux_stage_1[11] = (sel_1_reg0 == 1'b1) ? mux_stage_2[13] : mux_stage_2[11];
	assign mux_stage_1[12] = (sel_1_reg0 == 1'b1) ? mux_stage_2[14] : mux_stage_2[12];
	assign mux_stage_1[13] = (sel_1_reg0 == 1'b1) ? mux_stage_2[15] : mux_stage_2[13];
	assign mux_stage_1[14] = (sel_1_reg0 == 1'b1) ? mux_stage_2[16] : mux_stage_2[14];
	assign mux_stage_1[15] = (sel_1_reg0 == 1'b1) ? mux_stage_2[17] : mux_stage_2[15];
	assign mux_stage_1[16] = (sel_1_reg0 == 1'b1) ? mux_stage_2[18] : mux_stage_2[16];
	assign mux_stage_1[17] = (sel_1_reg0 == 1'b1) ? mux_stage_2[19] : mux_stage_2[17];
	assign mux_stage_1[18] = (sel_1_reg0 == 1'b1) ? mux_stage_2[20] : mux_stage_2[18];
	assign mux_stage_1[19] = (sel_1_reg0 == 1'b1) ? mux_stage_2[21] : mux_stage_2[19];
	assign mux_stage_1[20] = (sel_1_reg0 == 1'b1) ? mux_stage_2[22] : mux_stage_2[20];
	assign mux_stage_1[21] = (sel_1_reg0 == 1'b1) ? mux_stage_2[23] : mux_stage_2[21];
	assign mux_stage_1[22] = (sel_1_reg0 == 1'b1) ? mux_stage_2[24] : mux_stage_2[22];
	assign mux_stage_1[23] = (sel_1_reg0 == 1'b1) ? mux_stage_2[25] : mux_stage_2[23];
	assign mux_stage_1[24] = (sel_1_reg0 == 1'b1) ? mux_stage_2[26] : mux_stage_2[24];
	assign mux_stage_1[25] = (sel_1_reg0 == 1'b1) ? mux_stage_2[27] : mux_stage_2[25];
	assign mux_stage_1[26] = (sel_1_reg0 == 1'b1) ? mux_stage_2[28] : mux_stage_2[26];
	assign mux_stage_1[27] = (sel_1_reg0 == 1'b1) ? mux_stage_2[29] : mux_stage_2[27];
	assign mux_stage_1[28] = (sel_1_reg0 == 1'b1) ? mux_stage_2[30] : mux_stage_2[28];
	assign mux_stage_1[29] = (sel_1_reg0 == 1'b1) ? mux_stage_2[31] : mux_stage_2[29];
	assign mux_stage_1[30] = (sel_1_reg0 == 1'b1) ? mux_stage_2[32] : mux_stage_2[30];
	assign mux_stage_1[31] = (sel_1_reg0 == 1'b1) ? mux_stage_2[33] : mux_stage_2[31];
	assign mux_stage_1[32] = (sel_1_reg0 == 1'b1) ? mux_stage_2[34] : mux_stage_2[32];
	assign mux_stage_1[33] = (sel_1_reg0 == 1'b1) ? mux_stage_2[35] : mux_stage_2[33];
	assign mux_stage_1[34] = (sel_1_reg0 == 1'b1) ? mux_stage_2[36] : mux_stage_2[34];
	assign mux_stage_1[35] = (sel_1_reg0 == 1'b1) ? mux_stage_2[37] : mux_stage_2[35];
	assign mux_stage_1[36] = (sel_1_reg0 == 1'b1) ? mux_stage_2[38] : mux_stage_2[36];
	assign mux_stage_1[37] = (sel_1_reg0 == 1'b1) ? mux_stage_2[39] : mux_stage_2[37];
	assign mux_stage_1[38] = (sel_1_reg0 == 1'b1) ? mux_stage_2[40] : mux_stage_2[38];
	assign mux_stage_1[39] = (sel_1_reg0 == 1'b1) ? mux_stage_2[41] : mux_stage_2[39];
	assign mux_stage_1[40] = (sel_1_reg0 == 1'b1) ? mux_stage_2[42] : mux_stage_2[40];
	assign mux_stage_1[41] = (sel_1_reg0 == 1'b1) ? mux_stage_2[43] : mux_stage_2[41];
	assign mux_stage_1[42] = (sel_1_reg0 == 1'b1) ? mux_stage_2[44] : mux_stage_2[42];
	assign mux_stage_1[43] = (sel_1_reg0 == 1'b1) ? mux_stage_2[45] : mux_stage_2[43];
	assign mux_stage_1[44] = (sel_1_reg0 == 1'b1) ? mux_stage_2[46] : mux_stage_2[44];
	assign mux_stage_1[45] = (sel_1_reg0 == 1'b1) ? mux_stage_2[47] : mux_stage_2[45];
	assign mux_stage_1[46] = (sel_1_reg0 == 1'b1) ? mux_stage_2[48] : mux_stage_2[46];
	assign mux_stage_1[47] = (sel_1_reg0 == 1'b1) ? mux_stage_2[49] : mux_stage_2[47];
	assign mux_stage_1[48] = (sel_1_reg0 == 1'b1) ? mux_stage_2[50] : mux_stage_2[48];
	assign mux_stage_1[49] = (sel_1_reg0 == 1'b1) ? mux_stage_2[51] : mux_stage_2[49];
	assign mux_stage_1[50] = (sel_1_reg0 == 1'b1) ? mux_stage_2[52] : mux_stage_2[50];
	assign mux_stage_1[51] = (sel_1_reg0 == 1'b1) ? mux_stage_2[53] : mux_stage_2[51];
	assign mux_stage_1[52] = (sel_1_reg0 == 1'b1) ? mux_stage_2[54] : mux_stage_2[52];
	assign mux_stage_1[53] = (sel_1_reg0 == 1'b1) ? mux_stage_2[55] : mux_stage_2[53];
	assign mux_stage_1[54] = (sel_1_reg0 == 1'b1) ? mux_stage_2[56] : mux_stage_2[54];
	assign mux_stage_1[55] = (sel_1_reg0 == 1'b1) ? mux_stage_2[57] : mux_stage_2[55];
	assign mux_stage_1[56] = (sel_1_reg0 == 1'b1) ? mux_stage_2[58] : mux_stage_2[56];
	assign mux_stage_1[57] = (sel_1_reg0 == 1'b1) ? mux_stage_2[59] : mux_stage_2[57];
	assign mux_stage_1[58] = (sel_1_reg0 == 1'b1) ? mux_stage_2[60] : mux_stage_2[58];
	assign mux_stage_1[59] = (sel_1_reg0 == 1'b1) ? mux_stage_2[61] : mux_stage_2[59];
	assign mux_stage_1[60] = (sel_1_reg0 == 1'b1) ? mux_stage_2[62] : mux_stage_2[60];
	assign mux_stage_1[61] = (sel_1_reg0 == 1'b1) ? mux_stage_2[63] : mux_stage_2[61];
	assign mux_stage_1[62] = (sel_1_reg0 == 1'b1) ? mux_stage_2[64] : mux_stage_2[62];
	assign mux_stage_1[63] = (sel_1_reg0 == 1'b1) ? mux_stage_2[65] : mux_stage_2[63];
	assign mux_stage_1[64] = (sel_1_reg0 == 1'b1) ? mux_stage_2[66] : mux_stage_2[64];
	assign mux_stage_1[65] = (sel_1_reg0 == 1'b1) ? mux_stage_2[67] : mux_stage_2[65];
	assign mux_stage_1[66] = (sel_1_reg0 == 1'b1) ? mux_stage_2[68] : mux_stage_2[66];
	assign mux_stage_1[67] = (sel_1_reg0 == 1'b1) ? mux_stage_2[69] : mux_stage_2[67];
	assign mux_stage_1[68] = (sel_1_reg0 == 1'b1) ? mux_stage_2[70] : mux_stage_2[68];
	assign mux_stage_1[69] = (sel_1_reg0 == 1'b1) ? mux_stage_2[71] : mux_stage_2[69];
	assign mux_stage_1[70] = (sel_1_reg0 == 1'b1) ? mux_stage_2[72] : mux_stage_2[70];
	assign mux_stage_1[71] = (sel_1_reg0 == 1'b1) ? mux_stage_2[73] : mux_stage_2[71];
	assign mux_stage_1[72] = (sel_1_reg0 == 1'b1) ? mux_stage_2[74] : mux_stage_2[72];
	assign mux_stage_1[73] = (sel_1_reg0 == 1'b1) ? mux_stage_2[75] : mux_stage_2[73];
	assign mux_stage_1[74] = (sel_1_reg0 == 1'b1) ? mux_stage_2[76] : mux_stage_2[74];
	assign mux_stage_1[75] = (sel_1_reg0 == 1'b1) ? mux_stage_2[77] : mux_stage_2[75];
	assign mux_stage_1[76] = (sel_1_reg0 == 1'b1) ? mux_stage_2[78] : mux_stage_2[76];
	assign mux_stage_1[77] = (sel_1_reg0 == 1'b1) ? mux_stage_2[79] : mux_stage_2[77];
	assign mux_stage_1[78] = (sel_1_reg0 == 1'b1) ? mux_stage_2[80] : mux_stage_2[78];
	assign mux_stage_1[79] = (sel_1_reg0 == 1'b1) ? mux_stage_2[81] : mux_stage_2[79];
	assign mux_stage_1[80] = (sel_1_reg0 == 1'b1) ? mux_stage_2[82] : mux_stage_2[80];
	assign mux_stage_1[81] = (sel_1_reg0 == 1'b1) ? mux_stage_2[83] : mux_stage_2[81];
	assign mux_stage_1[82] = (sel_1_reg0 == 1'b1) ? mux_stage_2[84] : mux_stage_2[82];
	assign mux_stage_1[83] = (sel_1_reg0 == 1'b1) ? mux_stage_2[85] : mux_stage_2[83];
	assign mux_stage_1[84] = (sel_1_reg0 == 1'b1) ? mux_stage_2[86] : mux_stage_2[84];
	assign mux_stage_1[85] = (sel_1_reg0 == 1'b1) ? mux_stage_2[87] : mux_stage_2[85];
	assign mux_stage_1[86] = (sel_1_reg0 == 1'b1) ? mux_stage_2[88] : mux_stage_2[86];
	assign mux_stage_1[87] = (sel_1_reg0 == 1'b1) ? mux_stage_2[89] : mux_stage_2[87];
	assign mux_stage_1[88] = (sel_1_reg0 == 1'b1) ? mux_stage_2[90] : mux_stage_2[88];
	assign mux_stage_1[89] = (sel_1_reg0 == 1'b1) ? mux_stage_2[91] : mux_stage_2[89];
	assign mux_stage_1[90] = (sel_1_reg0 == 1'b1) ? mux_stage_2[92] : mux_stage_2[90];
	assign mux_stage_1[91] = (sel_1_reg0 == 1'b1) ? mux_stage_2[93] : mux_stage_2[91];
	assign mux_stage_1[92] = (sel_1_reg0 == 1'b1) ? mux_stage_2[94] : mux_stage_2[92];
	assign mux_stage_1[93] = (sel_1_reg0 == 1'b1) ? mux_stage_2[95] : mux_stage_2[93];
	assign mux_stage_1[94] = (sel_1_reg0 == 1'b1) ? mux_stage_2[96] : mux_stage_2[94];
	assign mux_stage_1[95] = (sel_1_reg0 == 1'b1) ? mux_stage_2[97] : mux_stage_2[95];
	assign mux_stage_1[96] = (sel_1_reg0 == 1'b1) ? mux_stage_2[98] : mux_stage_2[96];
	assign mux_stage_1[97] = (sel_1_reg0 == 1'b1) ? mux_stage_2[99] : mux_stage_2[97];
	assign mux_stage_1[98] = (sel_1_reg0 == 1'b1) ? mux_stage_2[100] : mux_stage_2[98];
	assign mux_stage_1[99] = (sel_1_reg0 == 1'b1) ? mux_stage_2[101] : mux_stage_2[99];
	assign mux_stage_1[100] = (sel_1_reg0 == 1'b1) ? mux_stage_2[102] : mux_stage_2[100];
	assign mux_stage_1[101] = (sel_1_reg0 == 1'b1) ? mux_stage_2[103] : mux_stage_2[101];
	assign mux_stage_1[102] = (sel_1_reg0 == 1'b1) ? mux_stage_2[104] : mux_stage_2[102];
	assign mux_stage_1[103] = (sel_1_reg0 == 1'b1) ? mux_stage_2[105] : mux_stage_2[103];
	assign mux_stage_1[104] = (sel_1_reg0 == 1'b1) ? mux_stage_2[106] : mux_stage_2[104];
	assign mux_stage_1[105] = (sel_1_reg0 == 1'b1) ? mux_stage_2[107] : mux_stage_2[105];
	assign mux_stage_1[106] = (sel_1_reg0 == 1'b1) ? mux_stage_2[108] : mux_stage_2[106];
	assign mux_stage_1[107] = (sel_1_reg0 == 1'b1) ? mux_stage_2[109] : mux_stage_2[107];
	assign mux_stage_1[108] = (sel_1_reg0 == 1'b1) ? mux_stage_2[110] : mux_stage_2[108];
	assign mux_stage_1[109] = (sel_1_reg0 == 1'b1) ? mux_stage_2[111] : mux_stage_2[109];
	assign mux_stage_1[110] = (sel_1_reg0 == 1'b1) ? mux_stage_2[112] : mux_stage_2[110];
	assign mux_stage_1[111] = (sel_1_reg0 == 1'b1) ? mux_stage_2[113] : mux_stage_2[111];
	assign mux_stage_1[112] = (sel_1_reg0 == 1'b1) ? mux_stage_2[114] : mux_stage_2[112];
	assign mux_stage_1[113] = (sel_1_reg0 == 1'b1) ? mux_stage_2[115] : mux_stage_2[113];
	assign mux_stage_1[114] = (sel_1_reg0 == 1'b1) ? mux_stage_2[116] : mux_stage_2[114];
	assign mux_stage_1[115] = (sel_1_reg0 == 1'b1) ? mux_stage_2[117] : mux_stage_2[115];
	assign mux_stage_1[116] = (sel_1_reg0 == 1'b1) ? mux_stage_2[118] : mux_stage_2[116];
	assign mux_stage_1[117] = (sel_1_reg0 == 1'b1) ? mux_stage_2[119] : mux_stage_2[117];
	assign mux_stage_1[118] = (sel_1_reg0 == 1'b1) ? mux_stage_2[120] : mux_stage_2[118];
	assign mux_stage_1[119] = (sel_1_reg0 == 1'b1) ? mux_stage_2[121] : mux_stage_2[119];
	assign mux_stage_1[120] = (sel_1_reg0 == 1'b1) ? mux_stage_2[122] : mux_stage_2[120];
	assign mux_stage_1[121] = (sel_1_reg0 == 1'b1) ? mux_stage_2[123] : mux_stage_2[121];
	assign mux_stage_1[122] = (sel_1_reg0 == 1'b1) ? mux_stage_2[124] : mux_stage_2[122];
	assign mux_stage_1[123] = (sel_1_reg0 == 1'b1) ? mux_stage_2[125] : mux_stage_2[123];
	assign mux_stage_1[124] = (sel_1_reg0 == 1'b1) ? mux_stage_2[126] : mux_stage_2[124];
	assign mux_stage_1[125] = (sel_1_reg0 == 1'b1) ? mux_stage_2[127] : mux_stage_2[125];
	assign mux_stage_1[126] = (sel_1_reg0 == 1'b1) ? mux_stage_2[128] : mux_stage_2[126];
	assign mux_stage_1[127] = (sel_1_reg0 == 1'b1) ? mux_stage_2[129] : mux_stage_2[127];
	assign mux_stage_1[128] = (sel_1_reg0 == 1'b1) ? mux_stage_2[130] : mux_stage_2[128];
	assign mux_stage_1[129] = (sel_1_reg0 == 1'b1) ? mux_stage_2[131] : mux_stage_2[129];
	assign mux_stage_1[130] = (sel_1_reg0 == 1'b1) ? mux_stage_2[132] : mux_stage_2[130];
	assign mux_stage_1[131] = (sel_1_reg0 == 1'b1) ? mux_stage_2[133] : mux_stage_2[131];
	assign mux_stage_1[132] = (sel_1_reg0 == 1'b1) ? mux_stage_2[134] : mux_stage_2[132];
	assign mux_stage_1[133] = (sel_1_reg0 == 1'b1) ? mux_stage_2[135] : mux_stage_2[133];
	assign mux_stage_1[134] = (sel_1_reg0 == 1'b1) ? mux_stage_2[136] : mux_stage_2[134];
	assign mux_stage_1[135] = (sel_1_reg0 == 1'b1) ? mux_stage_2[137] : mux_stage_2[135];
	assign mux_stage_1[136] = (sel_1_reg0 == 1'b1) ? mux_stage_2[138] : mux_stage_2[136];
	assign mux_stage_1[137] = (sel_1_reg0 == 1'b1) ? mux_stage_2[139] : mux_stage_2[137];
	assign mux_stage_1[138] = (sel_1_reg0 == 1'b1) ? mux_stage_2[140] : mux_stage_2[138];
	assign mux_stage_1[139] = (sel_1_reg0 == 1'b1) ? mux_stage_2[141] : mux_stage_2[139];
	assign mux_stage_1[140] = (sel_1_reg0 == 1'b1) ? mux_stage_2[142] : mux_stage_2[140];
	assign mux_stage_1[141] = (sel_1_reg0 == 1'b1) ? mux_stage_2[143] : mux_stage_2[141];
	assign mux_stage_1[142] = (sel_1_reg0 == 1'b1) ? mux_stage_2[144] : mux_stage_2[142];
	assign mux_stage_1[143] = (sel_1_reg0 == 1'b1) ? mux_stage_2[145] : mux_stage_2[143];
	assign mux_stage_1[144] = (sel_1_reg0 == 1'b1) ? mux_stage_2[146] : mux_stage_2[144];
	assign mux_stage_1[145] = (sel_1_reg0 == 1'b1) ? mux_stage_2[147] : mux_stage_2[145];
	assign mux_stage_1[146] = (sel_1_reg0 == 1'b1) ? mux_stage_2[148] : mux_stage_2[146];
	assign mux_stage_1[147] = (sel_1_reg0 == 1'b1) ? mux_stage_2[149] : mux_stage_2[147];
	assign mux_stage_1[148] = (sel_1_reg0 == 1'b1) ? mux_stage_2[150] : mux_stage_2[148];
	assign mux_stage_1[149] = (sel_1_reg0 == 1'b1) ? mux_stage_2[151] : mux_stage_2[149];
	assign mux_stage_1[150] = (sel_1_reg0 == 1'b1) ? mux_stage_2[152] : mux_stage_2[150];
	assign mux_stage_1[151] = (sel_1_reg0 == 1'b1) ? mux_stage_2[153] : mux_stage_2[151];
	assign mux_stage_1[152] = (sel_1_reg0 == 1'b1) ? mux_stage_2[154] : mux_stage_2[152];
	assign mux_stage_1[153] = (sel_1_reg0 == 1'b1) ? mux_stage_2[155] : mux_stage_2[153];
	assign mux_stage_1[154] = (sel_1_reg0 == 1'b1) ? mux_stage_2[156] : mux_stage_2[154];
	assign mux_stage_1[155] = (sel_1_reg0 == 1'b1) ? mux_stage_2[157] : mux_stage_2[155];
	assign mux_stage_1[156] = (sel_1_reg0 == 1'b1) ? mux_stage_2[158] : mux_stage_2[156];
	assign mux_stage_1[157] = (sel_1_reg0 == 1'b1) ? mux_stage_2[159] : mux_stage_2[157];
	assign mux_stage_1[158] = (sel_1_reg0 == 1'b1) ? mux_stage_2[160] : mux_stage_2[158];
	assign mux_stage_1[159] = (sel_1_reg0 == 1'b1) ? mux_stage_2[161] : mux_stage_2[159];
	assign mux_stage_1[160] = (sel_1_reg0 == 1'b1) ? mux_stage_2[162] : mux_stage_2[160];
	assign mux_stage_1[161] = (sel_1_reg0 == 1'b1) ? mux_stage_2[163] : mux_stage_2[161];
	assign mux_stage_1[162] = (sel_1_reg0 == 1'b1) ? mux_stage_2[164] : mux_stage_2[162];
	assign mux_stage_1[163] = (sel_1_reg0 == 1'b1) ? mux_stage_2[165] : mux_stage_2[163];
	assign mux_stage_1[164] = (sel_1_reg0 == 1'b1) ? mux_stage_2[166] : mux_stage_2[164];
	assign mux_stage_1[165] = (sel_1_reg0 == 1'b1) ? mux_stage_2[167] : mux_stage_2[165];
	assign mux_stage_1[166] = (sel_1_reg0 == 1'b1) ? mux_stage_2[168] : mux_stage_2[166];
	assign mux_stage_1[167] = (sel_1_reg0 == 1'b1) ? mux_stage_2[169] : mux_stage_2[167];
	assign mux_stage_1[168] = (sel_1_reg0 == 1'b1) ? mux_stage_2[170] : mux_stage_2[168];
	assign mux_stage_1[169] = (sel_1_reg0 == 1'b1) ? mux_stage_2[171] : mux_stage_2[169];
	assign mux_stage_1[170] = (sel_1_reg0 == 1'b1) ? mux_stage_2[172] : mux_stage_2[170];
	assign mux_stage_1[171] = (sel_1_reg0 == 1'b1) ? mux_stage_2[173] : mux_stage_2[171];
	assign mux_stage_1[172] = (sel_1_reg0 == 1'b1) ? mux_stage_2[174] : mux_stage_2[172];
	assign mux_stage_1[173] = (sel_1_reg0 == 1'b1) ? mux_stage_2[175] : mux_stage_2[173];
	assign mux_stage_1[174] = (sel_1_reg0 == 1'b1) ? mux_stage_2[176] : mux_stage_2[174];
	assign mux_stage_1[175] = (sel_1_reg0 == 1'b1) ? mux_stage_2[177] : mux_stage_2[175];
	assign mux_stage_1[176] = (sel_1_reg0 == 1'b1) ? mux_stage_2[178] : mux_stage_2[176];
	assign mux_stage_1[177] = (sel_1_reg0 == 1'b1) ? mux_stage_2[179] : mux_stage_2[177];
	assign mux_stage_1[178] = (sel_1_reg0 == 1'b1) ? mux_stage_2[180] : mux_stage_2[178];
	assign mux_stage_1[179] = (sel_1_reg0 == 1'b1) ? mux_stage_2[181] : mux_stage_2[179];
	assign mux_stage_1[180] = (sel_1_reg0 == 1'b1) ? mux_stage_2[182] : mux_stage_2[180];
	assign mux_stage_1[181] = (sel_1_reg0 == 1'b1) ? mux_stage_2[183] : mux_stage_2[181];
	assign mux_stage_1[182] = (sel_1_reg0 == 1'b1) ? mux_stage_2[184] : mux_stage_2[182];
	assign mux_stage_1[183] = (sel_1_reg0 == 1'b1) ? mux_stage_2[185] : mux_stage_2[183];
	assign mux_stage_1[184] = (sel_1_reg0 == 1'b1) ? mux_stage_2[186] : mux_stage_2[184];
	assign mux_stage_1[185] = (sel_1_reg0 == 1'b1) ? mux_stage_2[187] : mux_stage_2[185];
	assign mux_stage_1[186] = (sel_1_reg0 == 1'b1) ? mux_stage_2[188] : mux_stage_2[186];
	assign mux_stage_1[187] = (sel_1_reg0 == 1'b1) ? mux_stage_2[189] : mux_stage_2[187];
	assign mux_stage_1[188] = (sel_1_reg0 == 1'b1) ? mux_stage_2[190] : mux_stage_2[188];
	assign mux_stage_1[189] = (sel_1_reg0 == 1'b1) ? mux_stage_2[191] : mux_stage_2[189];
	assign mux_stage_1[190] = (sel_1_reg0 == 1'b1) ? mux_stage_2[192] : mux_stage_2[190];
	assign mux_stage_1[191] = (sel_1_reg0 == 1'b1) ? mux_stage_2[193] : mux_stage_2[191];
	assign mux_stage_1[192] = (sel_1_reg0 == 1'b1) ? mux_stage_2[194] : mux_stage_2[192];
	assign mux_stage_1[193] = (sel_1_reg0 == 1'b1) ? mux_stage_2[195] : mux_stage_2[193];
	assign mux_stage_1[194] = (sel_1_reg0 == 1'b1) ? mux_stage_2[196] : mux_stage_2[194];
	assign mux_stage_1[195] = (sel_1_reg0 == 1'b1) ? mux_stage_2[197] : mux_stage_2[195];
	assign mux_stage_1[196] = (sel_1_reg0 == 1'b1) ? mux_stage_2[198] : mux_stage_2[196];
	assign mux_stage_1[197] = (sel_1_reg0 == 1'b1) ? mux_stage_2[199] : mux_stage_2[197];
	assign mux_stage_1[198] = (sel_1_reg0 == 1'b1) ? mux_stage_2[200] : mux_stage_2[198];
	assign mux_stage_1[199] = (sel_1_reg0 == 1'b1) ? mux_stage_2[201] : mux_stage_2[199];
	assign mux_stage_1[200] = (sel_1_reg0 == 1'b1) ? mux_stage_2[202] : mux_stage_2[200];
	assign mux_stage_1[201] = (sel_1_reg0 == 1'b1) ? mux_stage_2[203] : mux_stage_2[201];
	assign mux_stage_1[202] = (sel_1_reg0 == 1'b1) ? mux_stage_2[204] : mux_stage_2[202];
	assign mux_stage_1[203] = (sel_1_reg0 == 1'b1) ? mux_stage_2[205] : mux_stage_2[203];
	assign mux_stage_1[204] = (sel_1_reg0 == 1'b1) ? mux_stage_2[206] : mux_stage_2[204];
	assign mux_stage_1[205] = (sel_1_reg0 == 1'b1) ? mux_stage_2[207] : mux_stage_2[205];
	assign mux_stage_1[206] = (sel_1_reg0 == 1'b1) ? mux_stage_2[208] : mux_stage_2[206];
	assign mux_stage_1[207] = (sel_1_reg0 == 1'b1) ? mux_stage_2[209] : mux_stage_2[207];
	assign mux_stage_1[208] = (sel_1_reg0 == 1'b1) ? mux_stage_2[210] : mux_stage_2[208];
	assign mux_stage_1[209] = (sel_1_reg0 == 1'b1) ? mux_stage_2[211] : mux_stage_2[209];
	assign mux_stage_1[210] = (sel_1_reg0 == 1'b1) ? mux_stage_2[212] : mux_stage_2[210];
	assign mux_stage_1[211] = (sel_1_reg0 == 1'b1) ? mux_stage_2[213] : mux_stage_2[211];
	assign mux_stage_1[212] = (sel_1_reg0 == 1'b1) ? mux_stage_2[214] : mux_stage_2[212];
	assign mux_stage_1[213] = (sel_1_reg0 == 1'b1) ? mux_stage_2[215] : mux_stage_2[213];
	assign mux_stage_1[214] = (sel_1_reg0 == 1'b1) ? mux_stage_2[216] : mux_stage_2[214];
	assign mux_stage_1[215] = (sel_1_reg0 == 1'b1) ? mux_stage_2[217] : mux_stage_2[215];
	assign mux_stage_1[216] = (sel_1_reg0 == 1'b1) ? mux_stage_2[218] : mux_stage_2[216];
	assign mux_stage_1[217] = (sel_1_reg0 == 1'b1) ? mux_stage_2[219] : mux_stage_2[217];
	assign mux_stage_1[218] = (sel_1_reg0 == 1'b1) ? mux_stage_2[220] : mux_stage_2[218];
	assign mux_stage_1[219] = (sel_1_reg0 == 1'b1) ? mux_stage_2[221] : mux_stage_2[219];
	assign mux_stage_1[220] = (sel_1_reg0 == 1'b1) ? mux_stage_2[222] : mux_stage_2[220];
	assign mux_stage_1[221] = (sel_1_reg0 == 1'b1) ? mux_stage_2[223] : mux_stage_2[221];
	assign mux_stage_1[222] = (sel_1_reg0 == 1'b1) ? mux_stage_2[224] : mux_stage_2[222];
	assign mux_stage_1[223] = (sel_1_reg0 == 1'b1) ? mux_stage_2[225] : mux_stage_2[223];
	assign mux_stage_1[224] = (sel_1_reg0 == 1'b1) ? mux_stage_2[226] : mux_stage_2[224];
	assign mux_stage_1[225] = (sel_1_reg0 == 1'b1) ? mux_stage_2[227] : mux_stage_2[225];
	assign mux_stage_1[226] = (sel_1_reg0 == 1'b1) ? mux_stage_2[228] : mux_stage_2[226];
	assign mux_stage_1[227] = (sel_1_reg0 == 1'b1) ? mux_stage_2[229] : mux_stage_2[227];
	assign mux_stage_1[228] = (sel_1_reg0 == 1'b1) ? mux_stage_2[230] : mux_stage_2[228];
	assign mux_stage_1[229] = (sel_1_reg0 == 1'b1) ? mux_stage_2[231] : mux_stage_2[229];
	assign mux_stage_1[230] = (sel_1_reg0 == 1'b1) ? mux_stage_2[232] : mux_stage_2[230];
	assign mux_stage_1[231] = (sel_1_reg0 == 1'b1) ? mux_stage_2[233] : mux_stage_2[231];
	assign mux_stage_1[232] = (sel_1_reg0 == 1'b1) ? mux_stage_2[234] : mux_stage_2[232];
	assign mux_stage_1[233] = (sel_1_reg0 == 1'b1) ? mux_stage_2[235] : mux_stage_2[233];
	assign mux_stage_1[234] = (sel_1_reg0 == 1'b1) ? mux_stage_2[236] : mux_stage_2[234];
	assign mux_stage_1[235] = (sel_1_reg0 == 1'b1) ? mux_stage_2[237] : mux_stage_2[235];
	assign mux_stage_1[236] = (sel_1_reg0 == 1'b1) ? mux_stage_2[238] : mux_stage_2[236];
	assign mux_stage_1[237] = (sel_1_reg0 == 1'b1) ? mux_stage_2[239] : mux_stage_2[237];
	assign mux_stage_1[238] = (sel_1_reg0 == 1'b1) ? mux_stage_2[240] : mux_stage_2[238];
	assign mux_stage_1[239] = (sel_1_reg0 == 1'b1) ? mux_stage_2[241] : mux_stage_2[239];
	assign mux_stage_1[240] = (sel_1_reg0 == 1'b1) ? mux_stage_2[242] : mux_stage_2[240];
	assign mux_stage_1[241] = (sel_1_reg0 == 1'b1) ? mux_stage_2[243] : mux_stage_2[241];
	assign mux_stage_1[242] = (sel_1_reg0 == 1'b1) ? mux_stage_2[244] : mux_stage_2[242];
	assign mux_stage_1[243] = (sel_1_reg0 == 1'b1) ? mux_stage_2[245] : mux_stage_2[243];
	assign mux_stage_1[244] = (sel_1_reg0 == 1'b1) ? mux_stage_2[246] : mux_stage_2[244];
	assign mux_stage_1[245] = (sel_1_reg0 == 1'b1) ? mux_stage_2[247] : mux_stage_2[245];
	assign mux_stage_1[246] = (sel_1_reg0 == 1'b1) ? mux_stage_2[248] : mux_stage_2[246];
	assign mux_stage_1[247] = (sel_1_reg0 == 1'b1) ? mux_stage_2[249] : mux_stage_2[247];
	assign mux_stage_1[248] = (sel_1_reg0 == 1'b1) ? mux_stage_2[250] : mux_stage_2[248];
	assign mux_stage_1[249] = (sel_1_reg0 == 1'b1) ? sw_in_251_reg0 : mux_stage_2[249];
	assign mux_stage_1[250] = (sel_1_reg0 == 1'b1) ? sw_in_252_reg0 : mux_stage_2[250];
	assign mux_stage_1[251] = (sel_1_reg0 == 1'b1) ? sw_in_253_reg0 : sw_in_251_reg0;
	assign mux_stage_1[252] = (sel_1_reg0 == 1'b1) ? sw_in_254_reg0 : sw_in_252_reg0;


	reg sel_0_reg0;
	always @(posedge sys_clk) begin if(!rstn) sel_0_reg0 <= 0; else sel_0_reg0 <= sel[0]; end	

	// Multiplexer Stage 0
	wire [253:0] mux_stage_0;
	assign mux_stage_0[0] = (sel_0_reg0 == 1'b1) ? mux_stage_1[1] : mux_stage_1[0];
	assign mux_stage_0[1] = (sel_0_reg0 == 1'b1) ? mux_stage_1[2] : mux_stage_1[1];
	assign mux_stage_0[2] = (sel_0_reg0 == 1'b1) ? mux_stage_1[3] : mux_stage_1[2];
	assign mux_stage_0[3] = (sel_0_reg0 == 1'b1) ? mux_stage_1[4] : mux_stage_1[3];
	assign mux_stage_0[4] = (sel_0_reg0 == 1'b1) ? mux_stage_1[5] : mux_stage_1[4];
	assign mux_stage_0[5] = (sel_0_reg0 == 1'b1) ? mux_stage_1[6] : mux_stage_1[5];
	assign mux_stage_0[6] = (sel_0_reg0 == 1'b1) ? mux_stage_1[7] : mux_stage_1[6];
	assign mux_stage_0[7] = (sel_0_reg0 == 1'b1) ? mux_stage_1[8] : mux_stage_1[7];
	assign mux_stage_0[8] = (sel_0_reg0 == 1'b1) ? mux_stage_1[9] : mux_stage_1[8];
	assign mux_stage_0[9] = (sel_0_reg0 == 1'b1) ? mux_stage_1[10] : mux_stage_1[9];
	assign mux_stage_0[10] = (sel_0_reg0 == 1'b1) ? mux_stage_1[11] : mux_stage_1[10];
	assign mux_stage_0[11] = (sel_0_reg0 == 1'b1) ? mux_stage_1[12] : mux_stage_1[11];
	assign mux_stage_0[12] = (sel_0_reg0 == 1'b1) ? mux_stage_1[13] : mux_stage_1[12];
	assign mux_stage_0[13] = (sel_0_reg0 == 1'b1) ? mux_stage_1[14] : mux_stage_1[13];
	assign mux_stage_0[14] = (sel_0_reg0 == 1'b1) ? mux_stage_1[15] : mux_stage_1[14];
	assign mux_stage_0[15] = (sel_0_reg0 == 1'b1) ? mux_stage_1[16] : mux_stage_1[15];
	assign mux_stage_0[16] = (sel_0_reg0 == 1'b1) ? mux_stage_1[17] : mux_stage_1[16];
	assign mux_stage_0[17] = (sel_0_reg0 == 1'b1) ? mux_stage_1[18] : mux_stage_1[17];
	assign mux_stage_0[18] = (sel_0_reg0 == 1'b1) ? mux_stage_1[19] : mux_stage_1[18];
	assign mux_stage_0[19] = (sel_0_reg0 == 1'b1) ? mux_stage_1[20] : mux_stage_1[19];
	assign mux_stage_0[20] = (sel_0_reg0 == 1'b1) ? mux_stage_1[21] : mux_stage_1[20];
	assign mux_stage_0[21] = (sel_0_reg0 == 1'b1) ? mux_stage_1[22] : mux_stage_1[21];
	assign mux_stage_0[22] = (sel_0_reg0 == 1'b1) ? mux_stage_1[23] : mux_stage_1[22];
	assign mux_stage_0[23] = (sel_0_reg0 == 1'b1) ? mux_stage_1[24] : mux_stage_1[23];
	assign mux_stage_0[24] = (sel_0_reg0 == 1'b1) ? mux_stage_1[25] : mux_stage_1[24];
	assign mux_stage_0[25] = (sel_0_reg0 == 1'b1) ? mux_stage_1[26] : mux_stage_1[25];
	assign mux_stage_0[26] = (sel_0_reg0 == 1'b1) ? mux_stage_1[27] : mux_stage_1[26];
	assign mux_stage_0[27] = (sel_0_reg0 == 1'b1) ? mux_stage_1[28] : mux_stage_1[27];
	assign mux_stage_0[28] = (sel_0_reg0 == 1'b1) ? mux_stage_1[29] : mux_stage_1[28];
	assign mux_stage_0[29] = (sel_0_reg0 == 1'b1) ? mux_stage_1[30] : mux_stage_1[29];
	assign mux_stage_0[30] = (sel_0_reg0 == 1'b1) ? mux_stage_1[31] : mux_stage_1[30];
	assign mux_stage_0[31] = (sel_0_reg0 == 1'b1) ? mux_stage_1[32] : mux_stage_1[31];
	assign mux_stage_0[32] = (sel_0_reg0 == 1'b1) ? mux_stage_1[33] : mux_stage_1[32];
	assign mux_stage_0[33] = (sel_0_reg0 == 1'b1) ? mux_stage_1[34] : mux_stage_1[33];
	assign mux_stage_0[34] = (sel_0_reg0 == 1'b1) ? mux_stage_1[35] : mux_stage_1[34];
	assign mux_stage_0[35] = (sel_0_reg0 == 1'b1) ? mux_stage_1[36] : mux_stage_1[35];
	assign mux_stage_0[36] = (sel_0_reg0 == 1'b1) ? mux_stage_1[37] : mux_stage_1[36];
	assign mux_stage_0[37] = (sel_0_reg0 == 1'b1) ? mux_stage_1[38] : mux_stage_1[37];
	assign mux_stage_0[38] = (sel_0_reg0 == 1'b1) ? mux_stage_1[39] : mux_stage_1[38];
	assign mux_stage_0[39] = (sel_0_reg0 == 1'b1) ? mux_stage_1[40] : mux_stage_1[39];
	assign mux_stage_0[40] = (sel_0_reg0 == 1'b1) ? mux_stage_1[41] : mux_stage_1[40];
	assign mux_stage_0[41] = (sel_0_reg0 == 1'b1) ? mux_stage_1[42] : mux_stage_1[41];
	assign mux_stage_0[42] = (sel_0_reg0 == 1'b1) ? mux_stage_1[43] : mux_stage_1[42];
	assign mux_stage_0[43] = (sel_0_reg0 == 1'b1) ? mux_stage_1[44] : mux_stage_1[43];
	assign mux_stage_0[44] = (sel_0_reg0 == 1'b1) ? mux_stage_1[45] : mux_stage_1[44];
	assign mux_stage_0[45] = (sel_0_reg0 == 1'b1) ? mux_stage_1[46] : mux_stage_1[45];
	assign mux_stage_0[46] = (sel_0_reg0 == 1'b1) ? mux_stage_1[47] : mux_stage_1[46];
	assign mux_stage_0[47] = (sel_0_reg0 == 1'b1) ? mux_stage_1[48] : mux_stage_1[47];
	assign mux_stage_0[48] = (sel_0_reg0 == 1'b1) ? mux_stage_1[49] : mux_stage_1[48];
	assign mux_stage_0[49] = (sel_0_reg0 == 1'b1) ? mux_stage_1[50] : mux_stage_1[49];
	assign mux_stage_0[50] = (sel_0_reg0 == 1'b1) ? mux_stage_1[51] : mux_stage_1[50];
	assign mux_stage_0[51] = (sel_0_reg0 == 1'b1) ? mux_stage_1[52] : mux_stage_1[51];
	assign mux_stage_0[52] = (sel_0_reg0 == 1'b1) ? mux_stage_1[53] : mux_stage_1[52];
	assign mux_stage_0[53] = (sel_0_reg0 == 1'b1) ? mux_stage_1[54] : mux_stage_1[53];
	assign mux_stage_0[54] = (sel_0_reg0 == 1'b1) ? mux_stage_1[55] : mux_stage_1[54];
	assign mux_stage_0[55] = (sel_0_reg0 == 1'b1) ? mux_stage_1[56] : mux_stage_1[55];
	assign mux_stage_0[56] = (sel_0_reg0 == 1'b1) ? mux_stage_1[57] : mux_stage_1[56];
	assign mux_stage_0[57] = (sel_0_reg0 == 1'b1) ? mux_stage_1[58] : mux_stage_1[57];
	assign mux_stage_0[58] = (sel_0_reg0 == 1'b1) ? mux_stage_1[59] : mux_stage_1[58];
	assign mux_stage_0[59] = (sel_0_reg0 == 1'b1) ? mux_stage_1[60] : mux_stage_1[59];
	assign mux_stage_0[60] = (sel_0_reg0 == 1'b1) ? mux_stage_1[61] : mux_stage_1[60];
	assign mux_stage_0[61] = (sel_0_reg0 == 1'b1) ? mux_stage_1[62] : mux_stage_1[61];
	assign mux_stage_0[62] = (sel_0_reg0 == 1'b1) ? mux_stage_1[63] : mux_stage_1[62];
	assign mux_stage_0[63] = (sel_0_reg0 == 1'b1) ? mux_stage_1[64] : mux_stage_1[63];
	assign mux_stage_0[64] = (sel_0_reg0 == 1'b1) ? mux_stage_1[65] : mux_stage_1[64];
	assign mux_stage_0[65] = (sel_0_reg0 == 1'b1) ? mux_stage_1[66] : mux_stage_1[65];
	assign mux_stage_0[66] = (sel_0_reg0 == 1'b1) ? mux_stage_1[67] : mux_stage_1[66];
	assign mux_stage_0[67] = (sel_0_reg0 == 1'b1) ? mux_stage_1[68] : mux_stage_1[67];
	assign mux_stage_0[68] = (sel_0_reg0 == 1'b1) ? mux_stage_1[69] : mux_stage_1[68];
	assign mux_stage_0[69] = (sel_0_reg0 == 1'b1) ? mux_stage_1[70] : mux_stage_1[69];
	assign mux_stage_0[70] = (sel_0_reg0 == 1'b1) ? mux_stage_1[71] : mux_stage_1[70];
	assign mux_stage_0[71] = (sel_0_reg0 == 1'b1) ? mux_stage_1[72] : mux_stage_1[71];
	assign mux_stage_0[72] = (sel_0_reg0 == 1'b1) ? mux_stage_1[73] : mux_stage_1[72];
	assign mux_stage_0[73] = (sel_0_reg0 == 1'b1) ? mux_stage_1[74] : mux_stage_1[73];
	assign mux_stage_0[74] = (sel_0_reg0 == 1'b1) ? mux_stage_1[75] : mux_stage_1[74];
	assign mux_stage_0[75] = (sel_0_reg0 == 1'b1) ? mux_stage_1[76] : mux_stage_1[75];
	assign mux_stage_0[76] = (sel_0_reg0 == 1'b1) ? mux_stage_1[77] : mux_stage_1[76];
	assign mux_stage_0[77] = (sel_0_reg0 == 1'b1) ? mux_stage_1[78] : mux_stage_1[77];
	assign mux_stage_0[78] = (sel_0_reg0 == 1'b1) ? mux_stage_1[79] : mux_stage_1[78];
	assign mux_stage_0[79] = (sel_0_reg0 == 1'b1) ? mux_stage_1[80] : mux_stage_1[79];
	assign mux_stage_0[80] = (sel_0_reg0 == 1'b1) ? mux_stage_1[81] : mux_stage_1[80];
	assign mux_stage_0[81] = (sel_0_reg0 == 1'b1) ? mux_stage_1[82] : mux_stage_1[81];
	assign mux_stage_0[82] = (sel_0_reg0 == 1'b1) ? mux_stage_1[83] : mux_stage_1[82];
	assign mux_stage_0[83] = (sel_0_reg0 == 1'b1) ? mux_stage_1[84] : mux_stage_1[83];
	assign mux_stage_0[84] = (sel_0_reg0 == 1'b1) ? mux_stage_1[85] : mux_stage_1[84];
	assign mux_stage_0[85] = (sel_0_reg0 == 1'b1) ? mux_stage_1[86] : mux_stage_1[85];
	assign mux_stage_0[86] = (sel_0_reg0 == 1'b1) ? mux_stage_1[87] : mux_stage_1[86];
	assign mux_stage_0[87] = (sel_0_reg0 == 1'b1) ? mux_stage_1[88] : mux_stage_1[87];
	assign mux_stage_0[88] = (sel_0_reg0 == 1'b1) ? mux_stage_1[89] : mux_stage_1[88];
	assign mux_stage_0[89] = (sel_0_reg0 == 1'b1) ? mux_stage_1[90] : mux_stage_1[89];
	assign mux_stage_0[90] = (sel_0_reg0 == 1'b1) ? mux_stage_1[91] : mux_stage_1[90];
	assign mux_stage_0[91] = (sel_0_reg0 == 1'b1) ? mux_stage_1[92] : mux_stage_1[91];
	assign mux_stage_0[92] = (sel_0_reg0 == 1'b1) ? mux_stage_1[93] : mux_stage_1[92];
	assign mux_stage_0[93] = (sel_0_reg0 == 1'b1) ? mux_stage_1[94] : mux_stage_1[93];
	assign mux_stage_0[94] = (sel_0_reg0 == 1'b1) ? mux_stage_1[95] : mux_stage_1[94];
	assign mux_stage_0[95] = (sel_0_reg0 == 1'b1) ? mux_stage_1[96] : mux_stage_1[95];
	assign mux_stage_0[96] = (sel_0_reg0 == 1'b1) ? mux_stage_1[97] : mux_stage_1[96];
	assign mux_stage_0[97] = (sel_0_reg0 == 1'b1) ? mux_stage_1[98] : mux_stage_1[97];
	assign mux_stage_0[98] = (sel_0_reg0 == 1'b1) ? mux_stage_1[99] : mux_stage_1[98];
	assign mux_stage_0[99] = (sel_0_reg0 == 1'b1) ? mux_stage_1[100] : mux_stage_1[99];
	assign mux_stage_0[100] = (sel_0_reg0 == 1'b1) ? mux_stage_1[101] : mux_stage_1[100];
	assign mux_stage_0[101] = (sel_0_reg0 == 1'b1) ? mux_stage_1[102] : mux_stage_1[101];
	assign mux_stage_0[102] = (sel_0_reg0 == 1'b1) ? mux_stage_1[103] : mux_stage_1[102];
	assign mux_stage_0[103] = (sel_0_reg0 == 1'b1) ? mux_stage_1[104] : mux_stage_1[103];
	assign mux_stage_0[104] = (sel_0_reg0 == 1'b1) ? mux_stage_1[105] : mux_stage_1[104];
	assign mux_stage_0[105] = (sel_0_reg0 == 1'b1) ? mux_stage_1[106] : mux_stage_1[105];
	assign mux_stage_0[106] = (sel_0_reg0 == 1'b1) ? mux_stage_1[107] : mux_stage_1[106];
	assign mux_stage_0[107] = (sel_0_reg0 == 1'b1) ? mux_stage_1[108] : mux_stage_1[107];
	assign mux_stage_0[108] = (sel_0_reg0 == 1'b1) ? mux_stage_1[109] : mux_stage_1[108];
	assign mux_stage_0[109] = (sel_0_reg0 == 1'b1) ? mux_stage_1[110] : mux_stage_1[109];
	assign mux_stage_0[110] = (sel_0_reg0 == 1'b1) ? mux_stage_1[111] : mux_stage_1[110];
	assign mux_stage_0[111] = (sel_0_reg0 == 1'b1) ? mux_stage_1[112] : mux_stage_1[111];
	assign mux_stage_0[112] = (sel_0_reg0 == 1'b1) ? mux_stage_1[113] : mux_stage_1[112];
	assign mux_stage_0[113] = (sel_0_reg0 == 1'b1) ? mux_stage_1[114] : mux_stage_1[113];
	assign mux_stage_0[114] = (sel_0_reg0 == 1'b1) ? mux_stage_1[115] : mux_stage_1[114];
	assign mux_stage_0[115] = (sel_0_reg0 == 1'b1) ? mux_stage_1[116] : mux_stage_1[115];
	assign mux_stage_0[116] = (sel_0_reg0 == 1'b1) ? mux_stage_1[117] : mux_stage_1[116];
	assign mux_stage_0[117] = (sel_0_reg0 == 1'b1) ? mux_stage_1[118] : mux_stage_1[117];
	assign mux_stage_0[118] = (sel_0_reg0 == 1'b1) ? mux_stage_1[119] : mux_stage_1[118];
	assign mux_stage_0[119] = (sel_0_reg0 == 1'b1) ? mux_stage_1[120] : mux_stage_1[119];
	assign mux_stage_0[120] = (sel_0_reg0 == 1'b1) ? mux_stage_1[121] : mux_stage_1[120];
	assign mux_stage_0[121] = (sel_0_reg0 == 1'b1) ? mux_stage_1[122] : mux_stage_1[121];
	assign mux_stage_0[122] = (sel_0_reg0 == 1'b1) ? mux_stage_1[123] : mux_stage_1[122];
	assign mux_stage_0[123] = (sel_0_reg0 == 1'b1) ? mux_stage_1[124] : mux_stage_1[123];
	assign mux_stage_0[124] = (sel_0_reg0 == 1'b1) ? mux_stage_1[125] : mux_stage_1[124];
	assign mux_stage_0[125] = (sel_0_reg0 == 1'b1) ? mux_stage_1[126] : mux_stage_1[125];
	assign mux_stage_0[126] = (sel_0_reg0 == 1'b1) ? mux_stage_1[127] : mux_stage_1[126];
	assign mux_stage_0[127] = (sel_0_reg0 == 1'b1) ? mux_stage_1[128] : mux_stage_1[127];
	assign mux_stage_0[128] = (sel_0_reg0 == 1'b1) ? mux_stage_1[129] : mux_stage_1[128];
	assign mux_stage_0[129] = (sel_0_reg0 == 1'b1) ? mux_stage_1[130] : mux_stage_1[129];
	assign mux_stage_0[130] = (sel_0_reg0 == 1'b1) ? mux_stage_1[131] : mux_stage_1[130];
	assign mux_stage_0[131] = (sel_0_reg0 == 1'b1) ? mux_stage_1[132] : mux_stage_1[131];
	assign mux_stage_0[132] = (sel_0_reg0 == 1'b1) ? mux_stage_1[133] : mux_stage_1[132];
	assign mux_stage_0[133] = (sel_0_reg0 == 1'b1) ? mux_stage_1[134] : mux_stage_1[133];
	assign mux_stage_0[134] = (sel_0_reg0 == 1'b1) ? mux_stage_1[135] : mux_stage_1[134];
	assign mux_stage_0[135] = (sel_0_reg0 == 1'b1) ? mux_stage_1[136] : mux_stage_1[135];
	assign mux_stage_0[136] = (sel_0_reg0 == 1'b1) ? mux_stage_1[137] : mux_stage_1[136];
	assign mux_stage_0[137] = (sel_0_reg0 == 1'b1) ? mux_stage_1[138] : mux_stage_1[137];
	assign mux_stage_0[138] = (sel_0_reg0 == 1'b1) ? mux_stage_1[139] : mux_stage_1[138];
	assign mux_stage_0[139] = (sel_0_reg0 == 1'b1) ? mux_stage_1[140] : mux_stage_1[139];
	assign mux_stage_0[140] = (sel_0_reg0 == 1'b1) ? mux_stage_1[141] : mux_stage_1[140];
	assign mux_stage_0[141] = (sel_0_reg0 == 1'b1) ? mux_stage_1[142] : mux_stage_1[141];
	assign mux_stage_0[142] = (sel_0_reg0 == 1'b1) ? mux_stage_1[143] : mux_stage_1[142];
	assign mux_stage_0[143] = (sel_0_reg0 == 1'b1) ? mux_stage_1[144] : mux_stage_1[143];
	assign mux_stage_0[144] = (sel_0_reg0 == 1'b1) ? mux_stage_1[145] : mux_stage_1[144];
	assign mux_stage_0[145] = (sel_0_reg0 == 1'b1) ? mux_stage_1[146] : mux_stage_1[145];
	assign mux_stage_0[146] = (sel_0_reg0 == 1'b1) ? mux_stage_1[147] : mux_stage_1[146];
	assign mux_stage_0[147] = (sel_0_reg0 == 1'b1) ? mux_stage_1[148] : mux_stage_1[147];
	assign mux_stage_0[148] = (sel_0_reg0 == 1'b1) ? mux_stage_1[149] : mux_stage_1[148];
	assign mux_stage_0[149] = (sel_0_reg0 == 1'b1) ? mux_stage_1[150] : mux_stage_1[149];
	assign mux_stage_0[150] = (sel_0_reg0 == 1'b1) ? mux_stage_1[151] : mux_stage_1[150];
	assign mux_stage_0[151] = (sel_0_reg0 == 1'b1) ? mux_stage_1[152] : mux_stage_1[151];
	assign mux_stage_0[152] = (sel_0_reg0 == 1'b1) ? mux_stage_1[153] : mux_stage_1[152];
	assign mux_stage_0[153] = (sel_0_reg0 == 1'b1) ? mux_stage_1[154] : mux_stage_1[153];
	assign mux_stage_0[154] = (sel_0_reg0 == 1'b1) ? mux_stage_1[155] : mux_stage_1[154];
	assign mux_stage_0[155] = (sel_0_reg0 == 1'b1) ? mux_stage_1[156] : mux_stage_1[155];
	assign mux_stage_0[156] = (sel_0_reg0 == 1'b1) ? mux_stage_1[157] : mux_stage_1[156];
	assign mux_stage_0[157] = (sel_0_reg0 == 1'b1) ? mux_stage_1[158] : mux_stage_1[157];
	assign mux_stage_0[158] = (sel_0_reg0 == 1'b1) ? mux_stage_1[159] : mux_stage_1[158];
	assign mux_stage_0[159] = (sel_0_reg0 == 1'b1) ? mux_stage_1[160] : mux_stage_1[159];
	assign mux_stage_0[160] = (sel_0_reg0 == 1'b1) ? mux_stage_1[161] : mux_stage_1[160];
	assign mux_stage_0[161] = (sel_0_reg0 == 1'b1) ? mux_stage_1[162] : mux_stage_1[161];
	assign mux_stage_0[162] = (sel_0_reg0 == 1'b1) ? mux_stage_1[163] : mux_stage_1[162];
	assign mux_stage_0[163] = (sel_0_reg0 == 1'b1) ? mux_stage_1[164] : mux_stage_1[163];
	assign mux_stage_0[164] = (sel_0_reg0 == 1'b1) ? mux_stage_1[165] : mux_stage_1[164];
	assign mux_stage_0[165] = (sel_0_reg0 == 1'b1) ? mux_stage_1[166] : mux_stage_1[165];
	assign mux_stage_0[166] = (sel_0_reg0 == 1'b1) ? mux_stage_1[167] : mux_stage_1[166];
	assign mux_stage_0[167] = (sel_0_reg0 == 1'b1) ? mux_stage_1[168] : mux_stage_1[167];
	assign mux_stage_0[168] = (sel_0_reg0 == 1'b1) ? mux_stage_1[169] : mux_stage_1[168];
	assign mux_stage_0[169] = (sel_0_reg0 == 1'b1) ? mux_stage_1[170] : mux_stage_1[169];
	assign mux_stage_0[170] = (sel_0_reg0 == 1'b1) ? mux_stage_1[171] : mux_stage_1[170];
	assign mux_stage_0[171] = (sel_0_reg0 == 1'b1) ? mux_stage_1[172] : mux_stage_1[171];
	assign mux_stage_0[172] = (sel_0_reg0 == 1'b1) ? mux_stage_1[173] : mux_stage_1[172];
	assign mux_stage_0[173] = (sel_0_reg0 == 1'b1) ? mux_stage_1[174] : mux_stage_1[173];
	assign mux_stage_0[174] = (sel_0_reg0 == 1'b1) ? mux_stage_1[175] : mux_stage_1[174];
	assign mux_stage_0[175] = (sel_0_reg0 == 1'b1) ? mux_stage_1[176] : mux_stage_1[175];
	assign mux_stage_0[176] = (sel_0_reg0 == 1'b1) ? mux_stage_1[177] : mux_stage_1[176];
	assign mux_stage_0[177] = (sel_0_reg0 == 1'b1) ? mux_stage_1[178] : mux_stage_1[177];
	assign mux_stage_0[178] = (sel_0_reg0 == 1'b1) ? mux_stage_1[179] : mux_stage_1[178];
	assign mux_stage_0[179] = (sel_0_reg0 == 1'b1) ? mux_stage_1[180] : mux_stage_1[179];
	assign mux_stage_0[180] = (sel_0_reg0 == 1'b1) ? mux_stage_1[181] : mux_stage_1[180];
	assign mux_stage_0[181] = (sel_0_reg0 == 1'b1) ? mux_stage_1[182] : mux_stage_1[181];
	assign mux_stage_0[182] = (sel_0_reg0 == 1'b1) ? mux_stage_1[183] : mux_stage_1[182];
	assign mux_stage_0[183] = (sel_0_reg0 == 1'b1) ? mux_stage_1[184] : mux_stage_1[183];
	assign mux_stage_0[184] = (sel_0_reg0 == 1'b1) ? mux_stage_1[185] : mux_stage_1[184];
	assign mux_stage_0[185] = (sel_0_reg0 == 1'b1) ? mux_stage_1[186] : mux_stage_1[185];
	assign mux_stage_0[186] = (sel_0_reg0 == 1'b1) ? mux_stage_1[187] : mux_stage_1[186];
	assign mux_stage_0[187] = (sel_0_reg0 == 1'b1) ? mux_stage_1[188] : mux_stage_1[187];
	assign mux_stage_0[188] = (sel_0_reg0 == 1'b1) ? mux_stage_1[189] : mux_stage_1[188];
	assign mux_stage_0[189] = (sel_0_reg0 == 1'b1) ? mux_stage_1[190] : mux_stage_1[189];
	assign mux_stage_0[190] = (sel_0_reg0 == 1'b1) ? mux_stage_1[191] : mux_stage_1[190];
	assign mux_stage_0[191] = (sel_0_reg0 == 1'b1) ? mux_stage_1[192] : mux_stage_1[191];
	assign mux_stage_0[192] = (sel_0_reg0 == 1'b1) ? mux_stage_1[193] : mux_stage_1[192];
	assign mux_stage_0[193] = (sel_0_reg0 == 1'b1) ? mux_stage_1[194] : mux_stage_1[193];
	assign mux_stage_0[194] = (sel_0_reg0 == 1'b1) ? mux_stage_1[195] : mux_stage_1[194];
	assign mux_stage_0[195] = (sel_0_reg0 == 1'b1) ? mux_stage_1[196] : mux_stage_1[195];
	assign mux_stage_0[196] = (sel_0_reg0 == 1'b1) ? mux_stage_1[197] : mux_stage_1[196];
	assign mux_stage_0[197] = (sel_0_reg0 == 1'b1) ? mux_stage_1[198] : mux_stage_1[197];
	assign mux_stage_0[198] = (sel_0_reg0 == 1'b1) ? mux_stage_1[199] : mux_stage_1[198];
	assign mux_stage_0[199] = (sel_0_reg0 == 1'b1) ? mux_stage_1[200] : mux_stage_1[199];
	assign mux_stage_0[200] = (sel_0_reg0 == 1'b1) ? mux_stage_1[201] : mux_stage_1[200];
	assign mux_stage_0[201] = (sel_0_reg0 == 1'b1) ? mux_stage_1[202] : mux_stage_1[201];
	assign mux_stage_0[202] = (sel_0_reg0 == 1'b1) ? mux_stage_1[203] : mux_stage_1[202];
	assign mux_stage_0[203] = (sel_0_reg0 == 1'b1) ? mux_stage_1[204] : mux_stage_1[203];
	assign mux_stage_0[204] = (sel_0_reg0 == 1'b1) ? mux_stage_1[205] : mux_stage_1[204];
	assign mux_stage_0[205] = (sel_0_reg0 == 1'b1) ? mux_stage_1[206] : mux_stage_1[205];
	assign mux_stage_0[206] = (sel_0_reg0 == 1'b1) ? mux_stage_1[207] : mux_stage_1[206];
	assign mux_stage_0[207] = (sel_0_reg0 == 1'b1) ? mux_stage_1[208] : mux_stage_1[207];
	assign mux_stage_0[208] = (sel_0_reg0 == 1'b1) ? mux_stage_1[209] : mux_stage_1[208];
	assign mux_stage_0[209] = (sel_0_reg0 == 1'b1) ? mux_stage_1[210] : mux_stage_1[209];
	assign mux_stage_0[210] = (sel_0_reg0 == 1'b1) ? mux_stage_1[211] : mux_stage_1[210];
	assign mux_stage_0[211] = (sel_0_reg0 == 1'b1) ? mux_stage_1[212] : mux_stage_1[211];
	assign mux_stage_0[212] = (sel_0_reg0 == 1'b1) ? mux_stage_1[213] : mux_stage_1[212];
	assign mux_stage_0[213] = (sel_0_reg0 == 1'b1) ? mux_stage_1[214] : mux_stage_1[213];
	assign mux_stage_0[214] = (sel_0_reg0 == 1'b1) ? mux_stage_1[215] : mux_stage_1[214];
	assign mux_stage_0[215] = (sel_0_reg0 == 1'b1) ? mux_stage_1[216] : mux_stage_1[215];
	assign mux_stage_0[216] = (sel_0_reg0 == 1'b1) ? mux_stage_1[217] : mux_stage_1[216];
	assign mux_stage_0[217] = (sel_0_reg0 == 1'b1) ? mux_stage_1[218] : mux_stage_1[217];
	assign mux_stage_0[218] = (sel_0_reg0 == 1'b1) ? mux_stage_1[219] : mux_stage_1[218];
	assign mux_stage_0[219] = (sel_0_reg0 == 1'b1) ? mux_stage_1[220] : mux_stage_1[219];
	assign mux_stage_0[220] = (sel_0_reg0 == 1'b1) ? mux_stage_1[221] : mux_stage_1[220];
	assign mux_stage_0[221] = (sel_0_reg0 == 1'b1) ? mux_stage_1[222] : mux_stage_1[221];
	assign mux_stage_0[222] = (sel_0_reg0 == 1'b1) ? mux_stage_1[223] : mux_stage_1[222];
	assign mux_stage_0[223] = (sel_0_reg0 == 1'b1) ? mux_stage_1[224] : mux_stage_1[223];
	assign mux_stage_0[224] = (sel_0_reg0 == 1'b1) ? mux_stage_1[225] : mux_stage_1[224];
	assign mux_stage_0[225] = (sel_0_reg0 == 1'b1) ? mux_stage_1[226] : mux_stage_1[225];
	assign mux_stage_0[226] = (sel_0_reg0 == 1'b1) ? mux_stage_1[227] : mux_stage_1[226];
	assign mux_stage_0[227] = (sel_0_reg0 == 1'b1) ? mux_stage_1[228] : mux_stage_1[227];
	assign mux_stage_0[228] = (sel_0_reg0 == 1'b1) ? mux_stage_1[229] : mux_stage_1[228];
	assign mux_stage_0[229] = (sel_0_reg0 == 1'b1) ? mux_stage_1[230] : mux_stage_1[229];
	assign mux_stage_0[230] = (sel_0_reg0 == 1'b1) ? mux_stage_1[231] : mux_stage_1[230];
	assign mux_stage_0[231] = (sel_0_reg0 == 1'b1) ? mux_stage_1[232] : mux_stage_1[231];
	assign mux_stage_0[232] = (sel_0_reg0 == 1'b1) ? mux_stage_1[233] : mux_stage_1[232];
	assign mux_stage_0[233] = (sel_0_reg0 == 1'b1) ? mux_stage_1[234] : mux_stage_1[233];
	assign mux_stage_0[234] = (sel_0_reg0 == 1'b1) ? mux_stage_1[235] : mux_stage_1[234];
	assign mux_stage_0[235] = (sel_0_reg0 == 1'b1) ? mux_stage_1[236] : mux_stage_1[235];
	assign mux_stage_0[236] = (sel_0_reg0 == 1'b1) ? mux_stage_1[237] : mux_stage_1[236];
	assign mux_stage_0[237] = (sel_0_reg0 == 1'b1) ? mux_stage_1[238] : mux_stage_1[237];
	assign mux_stage_0[238] = (sel_0_reg0 == 1'b1) ? mux_stage_1[239] : mux_stage_1[238];
	assign mux_stage_0[239] = (sel_0_reg0 == 1'b1) ? mux_stage_1[240] : mux_stage_1[239];
	assign mux_stage_0[240] = (sel_0_reg0 == 1'b1) ? mux_stage_1[241] : mux_stage_1[240];
	assign mux_stage_0[241] = (sel_0_reg0 == 1'b1) ? mux_stage_1[242] : mux_stage_1[241];
	assign mux_stage_0[242] = (sel_0_reg0 == 1'b1) ? mux_stage_1[243] : mux_stage_1[242];
	assign mux_stage_0[243] = (sel_0_reg0 == 1'b1) ? mux_stage_1[244] : mux_stage_1[243];
	assign mux_stage_0[244] = (sel_0_reg0 == 1'b1) ? mux_stage_1[245] : mux_stage_1[244];
	assign mux_stage_0[245] = (sel_0_reg0 == 1'b1) ? mux_stage_1[246] : mux_stage_1[245];
	assign mux_stage_0[246] = (sel_0_reg0 == 1'b1) ? mux_stage_1[247] : mux_stage_1[246];
	assign mux_stage_0[247] = (sel_0_reg0 == 1'b1) ? mux_stage_1[248] : mux_stage_1[247];
	assign mux_stage_0[248] = (sel_0_reg0 == 1'b1) ? mux_stage_1[249] : mux_stage_1[248];
	assign mux_stage_0[249] = (sel_0_reg0 == 1'b1) ? mux_stage_1[250] : mux_stage_1[249];
	assign mux_stage_0[250] = (sel_0_reg0 == 1'b1) ? mux_stage_1[251] : mux_stage_1[250];
	assign mux_stage_0[251] = (sel_0_reg0 == 1'b1) ? mux_stage_1[252] : mux_stage_1[251];
	assign mux_stage_0[252] = (sel_0_reg0 == 1'b1) ? sw_in_253_reg0 : mux_stage_1[252];
	assign mux_stage_0[253] = (sel_0_reg0 == 1'b1) ? sw_in_254_reg0 : sw_in_253_reg0;

	assign sw_out[253:0] = mux_stage_0[253:0];
endmodule