//`include "define.v"
`define QUAN_SIZE 4
`define IB_ADDR 8

module reconf_ib_lut (
	output reg [`QUAN_SIZE-1:0] t_c,
	
	input wire [`IB_ADDR-1:0] addr_in,
	input wire [`QUAN_SIZE-1:0] t_0,
	input wire [`QUAN_SIZE-1:0] t_1,
	input wire [`QUAN_SIZE-1:0] t_2,
	input wire [`QUAN_SIZE-1:0] t_3,
	input wire [`QUAN_SIZE-1:0] t_4,
	input wire [`QUAN_SIZE-1:0] t_5,
	input wire [`QUAN_SIZE-1:0] t_6,
	input wire [`QUAN_SIZE-1:0] t_7,
	input wire [`QUAN_SIZE-1:0] t_8,
	input wire [`QUAN_SIZE-1:0] t_9,
	input wire [`QUAN_SIZE-1:0] t_10,
	input wire [`QUAN_SIZE-1:0] t_11,
	input wire [`QUAN_SIZE-1:0] t_12,
	input wire [`QUAN_SIZE-1:0] t_13,
	input wire [`QUAN_SIZE-1:0] t_14,
	input wire [`QUAN_SIZE-1:0] t_15,
	input wire [`QUAN_SIZE-1:0] t_16,
	input wire [`QUAN_SIZE-1:0] t_17,
	input wire [`QUAN_SIZE-1:0] t_18,
	input wire [`QUAN_SIZE-1:0] t_19,
	input wire [`QUAN_SIZE-1:0] t_20,
	input wire [`QUAN_SIZE-1:0] t_21,
	input wire [`QUAN_SIZE-1:0] t_22,
	input wire [`QUAN_SIZE-1:0] t_23,
	input wire [`QUAN_SIZE-1:0] t_24,
	input wire [`QUAN_SIZE-1:0] t_25,
	input wire [`QUAN_SIZE-1:0] t_26,
	input wire [`QUAN_SIZE-1:0] t_27,
	input wire [`QUAN_SIZE-1:0] t_28,
	input wire [`QUAN_SIZE-1:0] t_29,
	input wire [`QUAN_SIZE-1:0] t_30,
	input wire [`QUAN_SIZE-1:0] t_31,
	input wire [`QUAN_SIZE-1:0] t_32,
	input wire [`QUAN_SIZE-1:0] t_33,
	input wire [`QUAN_SIZE-1:0] t_34,
	input wire [`QUAN_SIZE-1:0] t_35,
	input wire [`QUAN_SIZE-1:0] t_36,
	input wire [`QUAN_SIZE-1:0] t_37,
	input wire [`QUAN_SIZE-1:0] t_38,
	input wire [`QUAN_SIZE-1:0] t_39,
	input wire [`QUAN_SIZE-1:0] t_40,
	input wire [`QUAN_SIZE-1:0] t_41,
	input wire [`QUAN_SIZE-1:0] t_42,
	input wire [`QUAN_SIZE-1:0] t_43,
	input wire [`QUAN_SIZE-1:0] t_44,
	input wire [`QUAN_SIZE-1:0] t_45,
	input wire [`QUAN_SIZE-1:0] t_46,
	input wire [`QUAN_SIZE-1:0] t_47,
	input wire [`QUAN_SIZE-1:0] t_48,
	input wire [`QUAN_SIZE-1:0] t_49,
	input wire [`QUAN_SIZE-1:0] t_50,
	input wire [`QUAN_SIZE-1:0] t_51,
	input wire [`QUAN_SIZE-1:0] t_52,
	input wire [`QUAN_SIZE-1:0] t_53,
	input wire [`QUAN_SIZE-1:0] t_54,
	input wire [`QUAN_SIZE-1:0] t_55,
	input wire [`QUAN_SIZE-1:0] t_56,
	input wire [`QUAN_SIZE-1:0] t_57,
	input wire [`QUAN_SIZE-1:0] t_58,
	input wire [`QUAN_SIZE-1:0] t_59,
	input wire [`QUAN_SIZE-1:0] t_60,
	input wire [`QUAN_SIZE-1:0] t_61,
	input wire [`QUAN_SIZE-1:0] t_62,
	input wire [`QUAN_SIZE-1:0] t_63,
	input wire [`QUAN_SIZE-1:0] t_64,
	input wire [`QUAN_SIZE-1:0] t_65,
	input wire [`QUAN_SIZE-1:0] t_66,
	input wire [`QUAN_SIZE-1:0] t_67,
	input wire [`QUAN_SIZE-1:0] t_68,
	input wire [`QUAN_SIZE-1:0] t_69,
	input wire [`QUAN_SIZE-1:0] t_70,
	input wire [`QUAN_SIZE-1:0] t_71,
	input wire [`QUAN_SIZE-1:0] t_72,
	input wire [`QUAN_SIZE-1:0] t_73,
	input wire [`QUAN_SIZE-1:0] t_74,
	input wire [`QUAN_SIZE-1:0] t_75,
	input wire [`QUAN_SIZE-1:0] t_76,
	input wire [`QUAN_SIZE-1:0] t_77,
	input wire [`QUAN_SIZE-1:0] t_78,
	input wire [`QUAN_SIZE-1:0] t_79,
	input wire [`QUAN_SIZE-1:0] t_80,
	input wire [`QUAN_SIZE-1:0] t_81,
	input wire [`QUAN_SIZE-1:0] t_82,
	input wire [`QUAN_SIZE-1:0] t_83,
	input wire [`QUAN_SIZE-1:0] t_84,
	input wire [`QUAN_SIZE-1:0] t_85,
	input wire [`QUAN_SIZE-1:0] t_86,
	input wire [`QUAN_SIZE-1:0] t_87,
	input wire [`QUAN_SIZE-1:0] t_88,
	input wire [`QUAN_SIZE-1:0] t_89,
	input wire [`QUAN_SIZE-1:0] t_90,
	input wire [`QUAN_SIZE-1:0] t_91,
	input wire [`QUAN_SIZE-1:0] t_92,
	input wire [`QUAN_SIZE-1:0] t_93,
	input wire [`QUAN_SIZE-1:0] t_94,
	input wire [`QUAN_SIZE-1:0] t_95,
	input wire [`QUAN_SIZE-1:0] t_96,
	input wire [`QUAN_SIZE-1:0] t_97,
	input wire [`QUAN_SIZE-1:0] t_98,
	input wire [`QUAN_SIZE-1:0] t_99,
	input wire [`QUAN_SIZE-1:0] t_100,
	input wire [`QUAN_SIZE-1:0] t_101,
	input wire [`QUAN_SIZE-1:0] t_102,
	input wire [`QUAN_SIZE-1:0] t_103,
	input wire [`QUAN_SIZE-1:0] t_104,
	input wire [`QUAN_SIZE-1:0] t_105,
	input wire [`QUAN_SIZE-1:0] t_106,
	input wire [`QUAN_SIZE-1:0] t_107,
	input wire [`QUAN_SIZE-1:0] t_108,
	input wire [`QUAN_SIZE-1:0] t_109,
	input wire [`QUAN_SIZE-1:0] t_110,
	input wire [`QUAN_SIZE-1:0] t_111,
	input wire [`QUAN_SIZE-1:0] t_112,
	input wire [`QUAN_SIZE-1:0] t_113,
	input wire [`QUAN_SIZE-1:0] t_114,
	input wire [`QUAN_SIZE-1:0] t_115,
	input wire [`QUAN_SIZE-1:0] t_116,
	input wire [`QUAN_SIZE-1:0] t_117,
	input wire [`QUAN_SIZE-1:0] t_118,
	input wire [`QUAN_SIZE-1:0] t_119,
	input wire [`QUAN_SIZE-1:0] t_120,
	input wire [`QUAN_SIZE-1:0] t_121,
	input wire [`QUAN_SIZE-1:0] t_122,
	input wire [`QUAN_SIZE-1:0] t_123,
	input wire [`QUAN_SIZE-1:0] t_124,
	input wire [`QUAN_SIZE-1:0] t_125,
	input wire [`QUAN_SIZE-1:0] t_126,
	input wire [`QUAN_SIZE-1:0] t_127,
	input wire [`QUAN_SIZE-1:0] t_128,
	input wire [`QUAN_SIZE-1:0] t_129,
	input wire [`QUAN_SIZE-1:0] t_130,
	input wire [`QUAN_SIZE-1:0] t_131,
	input wire [`QUAN_SIZE-1:0] t_132,
	input wire [`QUAN_SIZE-1:0] t_133,
	input wire [`QUAN_SIZE-1:0] t_134,
	input wire [`QUAN_SIZE-1:0] t_135,
	input wire [`QUAN_SIZE-1:0] t_136,
	input wire [`QUAN_SIZE-1:0] t_137,
	input wire [`QUAN_SIZE-1:0] t_138,
	input wire [`QUAN_SIZE-1:0] t_139,
	input wire [`QUAN_SIZE-1:0] t_140,
	input wire [`QUAN_SIZE-1:0] t_141,
	input wire [`QUAN_SIZE-1:0] t_142,
	input wire [`QUAN_SIZE-1:0] t_143,
	input wire [`QUAN_SIZE-1:0] t_144,
	input wire [`QUAN_SIZE-1:0] t_145,
	input wire [`QUAN_SIZE-1:0] t_146,
	input wire [`QUAN_SIZE-1:0] t_147,
	input wire [`QUAN_SIZE-1:0] t_148,
	input wire [`QUAN_SIZE-1:0] t_149,
	input wire [`QUAN_SIZE-1:0] t_150,
	input wire [`QUAN_SIZE-1:0] t_151,
	input wire [`QUAN_SIZE-1:0] t_152,
	input wire [`QUAN_SIZE-1:0] t_153,
	input wire [`QUAN_SIZE-1:0] t_154,
	input wire [`QUAN_SIZE-1:0] t_155,
	input wire [`QUAN_SIZE-1:0] t_156,
	input wire [`QUAN_SIZE-1:0] t_157,
	input wire [`QUAN_SIZE-1:0] t_158,
	input wire [`QUAN_SIZE-1:0] t_159,
	input wire [`QUAN_SIZE-1:0] t_160,
	input wire [`QUAN_SIZE-1:0] t_161,
	input wire [`QUAN_SIZE-1:0] t_162,
	input wire [`QUAN_SIZE-1:0] t_163,
	input wire [`QUAN_SIZE-1:0] t_164,
	input wire [`QUAN_SIZE-1:0] t_165,
	input wire [`QUAN_SIZE-1:0] t_166,
	input wire [`QUAN_SIZE-1:0] t_167,
	input wire [`QUAN_SIZE-1:0] t_168,
	input wire [`QUAN_SIZE-1:0] t_169,
	input wire [`QUAN_SIZE-1:0] t_170,
	input wire [`QUAN_SIZE-1:0] t_171,
	input wire [`QUAN_SIZE-1:0] t_172,
	input wire [`QUAN_SIZE-1:0] t_173,
	input wire [`QUAN_SIZE-1:0] t_174,
	input wire [`QUAN_SIZE-1:0] t_175,
	input wire [`QUAN_SIZE-1:0] t_176,
	input wire [`QUAN_SIZE-1:0] t_177,
	input wire [`QUAN_SIZE-1:0] t_178,
	input wire [`QUAN_SIZE-1:0] t_179,
	input wire [`QUAN_SIZE-1:0] t_180,
	input wire [`QUAN_SIZE-1:0] t_181,
	input wire [`QUAN_SIZE-1:0] t_182,
	input wire [`QUAN_SIZE-1:0] t_183,
	input wire [`QUAN_SIZE-1:0] t_184,
	input wire [`QUAN_SIZE-1:0] t_185,
	input wire [`QUAN_SIZE-1:0] t_186,
	input wire [`QUAN_SIZE-1:0] t_187,
	input wire [`QUAN_SIZE-1:0] t_188,
	input wire [`QUAN_SIZE-1:0] t_189,
	input wire [`QUAN_SIZE-1:0] t_190,
	input wire [`QUAN_SIZE-1:0] t_191,
	input wire [`QUAN_SIZE-1:0] t_192,
	input wire [`QUAN_SIZE-1:0] t_193,
	input wire [`QUAN_SIZE-1:0] t_194,
	input wire [`QUAN_SIZE-1:0] t_195,
	input wire [`QUAN_SIZE-1:0] t_196,
	input wire [`QUAN_SIZE-1:0] t_197,
	input wire [`QUAN_SIZE-1:0] t_198,
	input wire [`QUAN_SIZE-1:0] t_199,
	input wire [`QUAN_SIZE-1:0] t_200,
	input wire [`QUAN_SIZE-1:0] t_201,
	input wire [`QUAN_SIZE-1:0] t_202,
	input wire [`QUAN_SIZE-1:0] t_203,
	input wire [`QUAN_SIZE-1:0] t_204,
	input wire [`QUAN_SIZE-1:0] t_205,
	input wire [`QUAN_SIZE-1:0] t_206,
	input wire [`QUAN_SIZE-1:0] t_207,
	input wire [`QUAN_SIZE-1:0] t_208,
	input wire [`QUAN_SIZE-1:0] t_209,
	input wire [`QUAN_SIZE-1:0] t_210,
	input wire [`QUAN_SIZE-1:0] t_211,
	input wire [`QUAN_SIZE-1:0] t_212,
	input wire [`QUAN_SIZE-1:0] t_213,
	input wire [`QUAN_SIZE-1:0] t_214,
	input wire [`QUAN_SIZE-1:0] t_215,
	input wire [`QUAN_SIZE-1:0] t_216,
	input wire [`QUAN_SIZE-1:0] t_217,
	input wire [`QUAN_SIZE-1:0] t_218,
	input wire [`QUAN_SIZE-1:0] t_219,
	input wire [`QUAN_SIZE-1:0] t_220,
	input wire [`QUAN_SIZE-1:0] t_221,
	input wire [`QUAN_SIZE-1:0] t_222,
	input wire [`QUAN_SIZE-1:0] t_223,
	input wire [`QUAN_SIZE-1:0] t_224,
	input wire [`QUAN_SIZE-1:0] t_225,
	input wire [`QUAN_SIZE-1:0] t_226,
	input wire [`QUAN_SIZE-1:0] t_227,
	input wire [`QUAN_SIZE-1:0] t_228,
	input wire [`QUAN_SIZE-1:0] t_229,
	input wire [`QUAN_SIZE-1:0] t_230,
	input wire [`QUAN_SIZE-1:0] t_231,
	input wire [`QUAN_SIZE-1:0] t_232,
	input wire [`QUAN_SIZE-1:0] t_233,
	input wire [`QUAN_SIZE-1:0] t_234,
	input wire [`QUAN_SIZE-1:0] t_235,
	input wire [`QUAN_SIZE-1:0] t_236,
	input wire [`QUAN_SIZE-1:0] t_237,
	input wire [`QUAN_SIZE-1:0] t_238,
	input wire [`QUAN_SIZE-1:0] t_239,
	input wire [`QUAN_SIZE-1:0] t_240,
	input wire [`QUAN_SIZE-1:0] t_241,
	input wire [`QUAN_SIZE-1:0] t_242,
	input wire [`QUAN_SIZE-1:0] t_243,
	input wire [`QUAN_SIZE-1:0] t_244,
	input wire [`QUAN_SIZE-1:0] t_245,
	input wire [`QUAN_SIZE-1:0] t_246,
	input wire [`QUAN_SIZE-1:0] t_247,
	input wire [`QUAN_SIZE-1:0] t_248,
	input wire [`QUAN_SIZE-1:0] t_249,
	input wire [`QUAN_SIZE-1:0] t_250,
	input wire [`QUAN_SIZE-1:0] t_251,
	input wire [`QUAN_SIZE-1:0] t_252,
	input wire [`QUAN_SIZE-1:0] t_253,
	input wire [`QUAN_SIZE-1:0] t_254,
	input wire [`QUAN_SIZE-1:0] t_255,

	input sys_clk
);

always @(posedge sys_clk) begin
	case(addr_in[`IB_ADDR-1:0])
		`IB_ADDR'd0: t_c[`QUAN_SIZE-1:0] = t_0[`QUAN_SIZE-1:0];
		`IB_ADDR'd1: t_c[`QUAN_SIZE-1:0] = t_1[`QUAN_SIZE-1:0];
		`IB_ADDR'd2: t_c[`QUAN_SIZE-1:0] = t_2[`QUAN_SIZE-1:0];
		`IB_ADDR'd3: t_c[`QUAN_SIZE-1:0] = t_3[`QUAN_SIZE-1:0];
		`IB_ADDR'd4: t_c[`QUAN_SIZE-1:0] = t_4[`QUAN_SIZE-1:0];
		`IB_ADDR'd5: t_c[`QUAN_SIZE-1:0] = t_5[`QUAN_SIZE-1:0];
		`IB_ADDR'd6: t_c[`QUAN_SIZE-1:0] = t_6[`QUAN_SIZE-1:0];
		`IB_ADDR'd7: t_c[`QUAN_SIZE-1:0] = t_7[`QUAN_SIZE-1:0];
		`IB_ADDR'd8: t_c[`QUAN_SIZE-1:0] = t_8[`QUAN_SIZE-1:0];
		`IB_ADDR'd9: t_c[`QUAN_SIZE-1:0] = t_9[`QUAN_SIZE-1:0];
		`IB_ADDR'd10: t_c[`QUAN_SIZE-1:0] = t_10[`QUAN_SIZE-1:0];
		`IB_ADDR'd11: t_c[`QUAN_SIZE-1:0] = t_11[`QUAN_SIZE-1:0];
		`IB_ADDR'd12: t_c[`QUAN_SIZE-1:0] = t_12[`QUAN_SIZE-1:0];
		`IB_ADDR'd13: t_c[`QUAN_SIZE-1:0] = t_13[`QUAN_SIZE-1:0];
		`IB_ADDR'd14: t_c[`QUAN_SIZE-1:0] = t_14[`QUAN_SIZE-1:0];
		`IB_ADDR'd15: t_c[`QUAN_SIZE-1:0] = t_15[`QUAN_SIZE-1:0];
		`IB_ADDR'd16: t_c[`QUAN_SIZE-1:0] = t_16[`QUAN_SIZE-1:0];
		`IB_ADDR'd17: t_c[`QUAN_SIZE-1:0] = t_17[`QUAN_SIZE-1:0];
		`IB_ADDR'd18: t_c[`QUAN_SIZE-1:0] = t_18[`QUAN_SIZE-1:0];
		`IB_ADDR'd19: t_c[`QUAN_SIZE-1:0] = t_19[`QUAN_SIZE-1:0];
		`IB_ADDR'd20: t_c[`QUAN_SIZE-1:0] = t_20[`QUAN_SIZE-1:0];
		`IB_ADDR'd21: t_c[`QUAN_SIZE-1:0] = t_21[`QUAN_SIZE-1:0];
		`IB_ADDR'd22: t_c[`QUAN_SIZE-1:0] = t_22[`QUAN_SIZE-1:0];
		`IB_ADDR'd23: t_c[`QUAN_SIZE-1:0] = t_23[`QUAN_SIZE-1:0];
		`IB_ADDR'd24: t_c[`QUAN_SIZE-1:0] = t_24[`QUAN_SIZE-1:0];
		`IB_ADDR'd25: t_c[`QUAN_SIZE-1:0] = t_25[`QUAN_SIZE-1:0];
		`IB_ADDR'd26: t_c[`QUAN_SIZE-1:0] = t_26[`QUAN_SIZE-1:0];
		`IB_ADDR'd27: t_c[`QUAN_SIZE-1:0] = t_27[`QUAN_SIZE-1:0];
		`IB_ADDR'd28: t_c[`QUAN_SIZE-1:0] = t_28[`QUAN_SIZE-1:0];
		`IB_ADDR'd29: t_c[`QUAN_SIZE-1:0] = t_29[`QUAN_SIZE-1:0];
		`IB_ADDR'd30: t_c[`QUAN_SIZE-1:0] = t_30[`QUAN_SIZE-1:0];
		`IB_ADDR'd31: t_c[`QUAN_SIZE-1:0] = t_31[`QUAN_SIZE-1:0];
		`IB_ADDR'd32: t_c[`QUAN_SIZE-1:0] = t_32[`QUAN_SIZE-1:0];
		`IB_ADDR'd33: t_c[`QUAN_SIZE-1:0] = t_33[`QUAN_SIZE-1:0];
		`IB_ADDR'd34: t_c[`QUAN_SIZE-1:0] = t_34[`QUAN_SIZE-1:0];
		`IB_ADDR'd35: t_c[`QUAN_SIZE-1:0] = t_35[`QUAN_SIZE-1:0];
		`IB_ADDR'd36: t_c[`QUAN_SIZE-1:0] = t_36[`QUAN_SIZE-1:0];
		`IB_ADDR'd37: t_c[`QUAN_SIZE-1:0] = t_37[`QUAN_SIZE-1:0];
		`IB_ADDR'd38: t_c[`QUAN_SIZE-1:0] = t_38[`QUAN_SIZE-1:0];
		`IB_ADDR'd39: t_c[`QUAN_SIZE-1:0] = t_39[`QUAN_SIZE-1:0];
		`IB_ADDR'd40: t_c[`QUAN_SIZE-1:0] = t_40[`QUAN_SIZE-1:0];
		`IB_ADDR'd41: t_c[`QUAN_SIZE-1:0] = t_41[`QUAN_SIZE-1:0];
		`IB_ADDR'd42: t_c[`QUAN_SIZE-1:0] = t_42[`QUAN_SIZE-1:0];
		`IB_ADDR'd43: t_c[`QUAN_SIZE-1:0] = t_43[`QUAN_SIZE-1:0];
		`IB_ADDR'd44: t_c[`QUAN_SIZE-1:0] = t_44[`QUAN_SIZE-1:0];
		`IB_ADDR'd45: t_c[`QUAN_SIZE-1:0] = t_45[`QUAN_SIZE-1:0];
		`IB_ADDR'd46: t_c[`QUAN_SIZE-1:0] = t_46[`QUAN_SIZE-1:0];
		`IB_ADDR'd47: t_c[`QUAN_SIZE-1:0] = t_47[`QUAN_SIZE-1:0];
		`IB_ADDR'd48: t_c[`QUAN_SIZE-1:0] = t_48[`QUAN_SIZE-1:0];
		`IB_ADDR'd49: t_c[`QUAN_SIZE-1:0] = t_49[`QUAN_SIZE-1:0];
		`IB_ADDR'd50: t_c[`QUAN_SIZE-1:0] = t_50[`QUAN_SIZE-1:0];
		`IB_ADDR'd51: t_c[`QUAN_SIZE-1:0] = t_51[`QUAN_SIZE-1:0];
		`IB_ADDR'd52: t_c[`QUAN_SIZE-1:0] = t_52[`QUAN_SIZE-1:0];
		`IB_ADDR'd53: t_c[`QUAN_SIZE-1:0] = t_53[`QUAN_SIZE-1:0];
		`IB_ADDR'd54: t_c[`QUAN_SIZE-1:0] = t_54[`QUAN_SIZE-1:0];
		`IB_ADDR'd55: t_c[`QUAN_SIZE-1:0] = t_55[`QUAN_SIZE-1:0];
		`IB_ADDR'd56: t_c[`QUAN_SIZE-1:0] = t_56[`QUAN_SIZE-1:0];
		`IB_ADDR'd57: t_c[`QUAN_SIZE-1:0] = t_57[`QUAN_SIZE-1:0];
		`IB_ADDR'd58: t_c[`QUAN_SIZE-1:0] = t_58[`QUAN_SIZE-1:0];
		`IB_ADDR'd59: t_c[`QUAN_SIZE-1:0] = t_59[`QUAN_SIZE-1:0];
		`IB_ADDR'd60: t_c[`QUAN_SIZE-1:0] = t_60[`QUAN_SIZE-1:0];
		`IB_ADDR'd61: t_c[`QUAN_SIZE-1:0] = t_61[`QUAN_SIZE-1:0];
		`IB_ADDR'd62: t_c[`QUAN_SIZE-1:0] = t_62[`QUAN_SIZE-1:0];
		`IB_ADDR'd63: t_c[`QUAN_SIZE-1:0] = t_63[`QUAN_SIZE-1:0];
		`IB_ADDR'd64: t_c[`QUAN_SIZE-1:0] = t_64[`QUAN_SIZE-1:0];
		`IB_ADDR'd65: t_c[`QUAN_SIZE-1:0] = t_65[`QUAN_SIZE-1:0];
		`IB_ADDR'd66: t_c[`QUAN_SIZE-1:0] = t_66[`QUAN_SIZE-1:0];
		`IB_ADDR'd67: t_c[`QUAN_SIZE-1:0] = t_67[`QUAN_SIZE-1:0];
		`IB_ADDR'd68: t_c[`QUAN_SIZE-1:0] = t_68[`QUAN_SIZE-1:0];
		`IB_ADDR'd69: t_c[`QUAN_SIZE-1:0] = t_69[`QUAN_SIZE-1:0];
		`IB_ADDR'd70: t_c[`QUAN_SIZE-1:0] = t_70[`QUAN_SIZE-1:0];
		`IB_ADDR'd71: t_c[`QUAN_SIZE-1:0] = t_71[`QUAN_SIZE-1:0];
		`IB_ADDR'd72: t_c[`QUAN_SIZE-1:0] = t_72[`QUAN_SIZE-1:0];
		`IB_ADDR'd73: t_c[`QUAN_SIZE-1:0] = t_73[`QUAN_SIZE-1:0];
		`IB_ADDR'd74: t_c[`QUAN_SIZE-1:0] = t_74[`QUAN_SIZE-1:0];
		`IB_ADDR'd75: t_c[`QUAN_SIZE-1:0] = t_75[`QUAN_SIZE-1:0];
		`IB_ADDR'd76: t_c[`QUAN_SIZE-1:0] = t_76[`QUAN_SIZE-1:0];
		`IB_ADDR'd77: t_c[`QUAN_SIZE-1:0] = t_77[`QUAN_SIZE-1:0];
		`IB_ADDR'd78: t_c[`QUAN_SIZE-1:0] = t_78[`QUAN_SIZE-1:0];
		`IB_ADDR'd79: t_c[`QUAN_SIZE-1:0] = t_79[`QUAN_SIZE-1:0];
		`IB_ADDR'd80: t_c[`QUAN_SIZE-1:0] = t_80[`QUAN_SIZE-1:0];
		`IB_ADDR'd81: t_c[`QUAN_SIZE-1:0] = t_81[`QUAN_SIZE-1:0];
		`IB_ADDR'd82: t_c[`QUAN_SIZE-1:0] = t_82[`QUAN_SIZE-1:0];
		`IB_ADDR'd83: t_c[`QUAN_SIZE-1:0] = t_83[`QUAN_SIZE-1:0];
		`IB_ADDR'd84: t_c[`QUAN_SIZE-1:0] = t_84[`QUAN_SIZE-1:0];
		`IB_ADDR'd85: t_c[`QUAN_SIZE-1:0] = t_85[`QUAN_SIZE-1:0];
		`IB_ADDR'd86: t_c[`QUAN_SIZE-1:0] = t_86[`QUAN_SIZE-1:0];
		`IB_ADDR'd87: t_c[`QUAN_SIZE-1:0] = t_87[`QUAN_SIZE-1:0];
		`IB_ADDR'd88: t_c[`QUAN_SIZE-1:0] = t_88[`QUAN_SIZE-1:0];
		`IB_ADDR'd89: t_c[`QUAN_SIZE-1:0] = t_89[`QUAN_SIZE-1:0];
		`IB_ADDR'd90: t_c[`QUAN_SIZE-1:0] = t_90[`QUAN_SIZE-1:0];
		`IB_ADDR'd91: t_c[`QUAN_SIZE-1:0] = t_91[`QUAN_SIZE-1:0];
		`IB_ADDR'd92: t_c[`QUAN_SIZE-1:0] = t_92[`QUAN_SIZE-1:0];
		`IB_ADDR'd93: t_c[`QUAN_SIZE-1:0] = t_93[`QUAN_SIZE-1:0];
		`IB_ADDR'd94: t_c[`QUAN_SIZE-1:0] = t_94[`QUAN_SIZE-1:0];
		`IB_ADDR'd95: t_c[`QUAN_SIZE-1:0] = t_95[`QUAN_SIZE-1:0];
		`IB_ADDR'd96: t_c[`QUAN_SIZE-1:0] = t_96[`QUAN_SIZE-1:0];
		`IB_ADDR'd97: t_c[`QUAN_SIZE-1:0] = t_97[`QUAN_SIZE-1:0];
		`IB_ADDR'd98: t_c[`QUAN_SIZE-1:0] = t_98[`QUAN_SIZE-1:0];
		`IB_ADDR'd99: t_c[`QUAN_SIZE-1:0] = t_99[`QUAN_SIZE-1:0];
		`IB_ADDR'd100: t_c[`QUAN_SIZE-1:0] = t_100[`QUAN_SIZE-1:0];
		`IB_ADDR'd101: t_c[`QUAN_SIZE-1:0] = t_101[`QUAN_SIZE-1:0];
		`IB_ADDR'd102: t_c[`QUAN_SIZE-1:0] = t_102[`QUAN_SIZE-1:0];
		`IB_ADDR'd103: t_c[`QUAN_SIZE-1:0] = t_103[`QUAN_SIZE-1:0];
		`IB_ADDR'd104: t_c[`QUAN_SIZE-1:0] = t_104[`QUAN_SIZE-1:0];
		`IB_ADDR'd105: t_c[`QUAN_SIZE-1:0] = t_105[`QUAN_SIZE-1:0];
		`IB_ADDR'd106: t_c[`QUAN_SIZE-1:0] = t_106[`QUAN_SIZE-1:0];
		`IB_ADDR'd107: t_c[`QUAN_SIZE-1:0] = t_107[`QUAN_SIZE-1:0];
		`IB_ADDR'd108: t_c[`QUAN_SIZE-1:0] = t_108[`QUAN_SIZE-1:0];
		`IB_ADDR'd109: t_c[`QUAN_SIZE-1:0] = t_109[`QUAN_SIZE-1:0];
		`IB_ADDR'd110: t_c[`QUAN_SIZE-1:0] = t_110[`QUAN_SIZE-1:0];
		`IB_ADDR'd111: t_c[`QUAN_SIZE-1:0] = t_111[`QUAN_SIZE-1:0];
		`IB_ADDR'd112: t_c[`QUAN_SIZE-1:0] = t_112[`QUAN_SIZE-1:0];
		`IB_ADDR'd113: t_c[`QUAN_SIZE-1:0] = t_113[`QUAN_SIZE-1:0];
		`IB_ADDR'd114: t_c[`QUAN_SIZE-1:0] = t_114[`QUAN_SIZE-1:0];
		`IB_ADDR'd115: t_c[`QUAN_SIZE-1:0] = t_115[`QUAN_SIZE-1:0];
		`IB_ADDR'd116: t_c[`QUAN_SIZE-1:0] = t_116[`QUAN_SIZE-1:0];
		`IB_ADDR'd117: t_c[`QUAN_SIZE-1:0] = t_117[`QUAN_SIZE-1:0];
		`IB_ADDR'd118: t_c[`QUAN_SIZE-1:0] = t_118[`QUAN_SIZE-1:0];
		`IB_ADDR'd119: t_c[`QUAN_SIZE-1:0] = t_119[`QUAN_SIZE-1:0];
		`IB_ADDR'd120: t_c[`QUAN_SIZE-1:0] = t_120[`QUAN_SIZE-1:0];
		`IB_ADDR'd121: t_c[`QUAN_SIZE-1:0] = t_121[`QUAN_SIZE-1:0];
		`IB_ADDR'd122: t_c[`QUAN_SIZE-1:0] = t_122[`QUAN_SIZE-1:0];
		`IB_ADDR'd123: t_c[`QUAN_SIZE-1:0] = t_123[`QUAN_SIZE-1:0];
		`IB_ADDR'd124: t_c[`QUAN_SIZE-1:0] = t_124[`QUAN_SIZE-1:0];
		`IB_ADDR'd125: t_c[`QUAN_SIZE-1:0] = t_125[`QUAN_SIZE-1:0];
		`IB_ADDR'd126: t_c[`QUAN_SIZE-1:0] = t_126[`QUAN_SIZE-1:0];
		`IB_ADDR'd127: t_c[`QUAN_SIZE-1:0] = t_127[`QUAN_SIZE-1:0];
		`IB_ADDR'd128: t_c[`QUAN_SIZE-1:0] = t_128[`QUAN_SIZE-1:0];
		`IB_ADDR'd129: t_c[`QUAN_SIZE-1:0] = t_129[`QUAN_SIZE-1:0];
		`IB_ADDR'd130: t_c[`QUAN_SIZE-1:0] = t_130[`QUAN_SIZE-1:0];
		`IB_ADDR'd131: t_c[`QUAN_SIZE-1:0] = t_131[`QUAN_SIZE-1:0];
		`IB_ADDR'd132: t_c[`QUAN_SIZE-1:0] = t_132[`QUAN_SIZE-1:0];
		`IB_ADDR'd133: t_c[`QUAN_SIZE-1:0] = t_133[`QUAN_SIZE-1:0];
		`IB_ADDR'd134: t_c[`QUAN_SIZE-1:0] = t_134[`QUAN_SIZE-1:0];
		`IB_ADDR'd135: t_c[`QUAN_SIZE-1:0] = t_135[`QUAN_SIZE-1:0];
		`IB_ADDR'd136: t_c[`QUAN_SIZE-1:0] = t_136[`QUAN_SIZE-1:0];
		`IB_ADDR'd137: t_c[`QUAN_SIZE-1:0] = t_137[`QUAN_SIZE-1:0];
		`IB_ADDR'd138: t_c[`QUAN_SIZE-1:0] = t_138[`QUAN_SIZE-1:0];
		`IB_ADDR'd139: t_c[`QUAN_SIZE-1:0] = t_139[`QUAN_SIZE-1:0];
		`IB_ADDR'd140: t_c[`QUAN_SIZE-1:0] = t_140[`QUAN_SIZE-1:0];
		`IB_ADDR'd141: t_c[`QUAN_SIZE-1:0] = t_141[`QUAN_SIZE-1:0];
		`IB_ADDR'd142: t_c[`QUAN_SIZE-1:0] = t_142[`QUAN_SIZE-1:0];
		`IB_ADDR'd143: t_c[`QUAN_SIZE-1:0] = t_143[`QUAN_SIZE-1:0];
		`IB_ADDR'd144: t_c[`QUAN_SIZE-1:0] = t_144[`QUAN_SIZE-1:0];
		`IB_ADDR'd145: t_c[`QUAN_SIZE-1:0] = t_145[`QUAN_SIZE-1:0];
		`IB_ADDR'd146: t_c[`QUAN_SIZE-1:0] = t_146[`QUAN_SIZE-1:0];
		`IB_ADDR'd147: t_c[`QUAN_SIZE-1:0] = t_147[`QUAN_SIZE-1:0];
		`IB_ADDR'd148: t_c[`QUAN_SIZE-1:0] = t_148[`QUAN_SIZE-1:0];
		`IB_ADDR'd149: t_c[`QUAN_SIZE-1:0] = t_149[`QUAN_SIZE-1:0];
		`IB_ADDR'd150: t_c[`QUAN_SIZE-1:0] = t_150[`QUAN_SIZE-1:0];
		`IB_ADDR'd151: t_c[`QUAN_SIZE-1:0] = t_151[`QUAN_SIZE-1:0];
		`IB_ADDR'd152: t_c[`QUAN_SIZE-1:0] = t_152[`QUAN_SIZE-1:0];
		`IB_ADDR'd153: t_c[`QUAN_SIZE-1:0] = t_153[`QUAN_SIZE-1:0];
		`IB_ADDR'd154: t_c[`QUAN_SIZE-1:0] = t_154[`QUAN_SIZE-1:0];
		`IB_ADDR'd155: t_c[`QUAN_SIZE-1:0] = t_155[`QUAN_SIZE-1:0];
		`IB_ADDR'd156: t_c[`QUAN_SIZE-1:0] = t_156[`QUAN_SIZE-1:0];
		`IB_ADDR'd157: t_c[`QUAN_SIZE-1:0] = t_157[`QUAN_SIZE-1:0];
		`IB_ADDR'd158: t_c[`QUAN_SIZE-1:0] = t_158[`QUAN_SIZE-1:0];
		`IB_ADDR'd159: t_c[`QUAN_SIZE-1:0] = t_159[`QUAN_SIZE-1:0];
		`IB_ADDR'd160: t_c[`QUAN_SIZE-1:0] = t_160[`QUAN_SIZE-1:0];
		`IB_ADDR'd161: t_c[`QUAN_SIZE-1:0] = t_161[`QUAN_SIZE-1:0];
		`IB_ADDR'd162: t_c[`QUAN_SIZE-1:0] = t_162[`QUAN_SIZE-1:0];
		`IB_ADDR'd163: t_c[`QUAN_SIZE-1:0] = t_163[`QUAN_SIZE-1:0];
		`IB_ADDR'd164: t_c[`QUAN_SIZE-1:0] = t_164[`QUAN_SIZE-1:0];
		`IB_ADDR'd165: t_c[`QUAN_SIZE-1:0] = t_165[`QUAN_SIZE-1:0];
		`IB_ADDR'd166: t_c[`QUAN_SIZE-1:0] = t_166[`QUAN_SIZE-1:0];
		`IB_ADDR'd167: t_c[`QUAN_SIZE-1:0] = t_167[`QUAN_SIZE-1:0];
		`IB_ADDR'd168: t_c[`QUAN_SIZE-1:0] = t_168[`QUAN_SIZE-1:0];
		`IB_ADDR'd169: t_c[`QUAN_SIZE-1:0] = t_169[`QUAN_SIZE-1:0];
		`IB_ADDR'd170: t_c[`QUAN_SIZE-1:0] = t_170[`QUAN_SIZE-1:0];
		`IB_ADDR'd171: t_c[`QUAN_SIZE-1:0] = t_171[`QUAN_SIZE-1:0];
		`IB_ADDR'd172: t_c[`QUAN_SIZE-1:0] = t_172[`QUAN_SIZE-1:0];
		`IB_ADDR'd173: t_c[`QUAN_SIZE-1:0] = t_173[`QUAN_SIZE-1:0];
		`IB_ADDR'd174: t_c[`QUAN_SIZE-1:0] = t_174[`QUAN_SIZE-1:0];
		`IB_ADDR'd175: t_c[`QUAN_SIZE-1:0] = t_175[`QUAN_SIZE-1:0];
		`IB_ADDR'd176: t_c[`QUAN_SIZE-1:0] = t_176[`QUAN_SIZE-1:0];
		`IB_ADDR'd177: t_c[`QUAN_SIZE-1:0] = t_177[`QUAN_SIZE-1:0];
		`IB_ADDR'd178: t_c[`QUAN_SIZE-1:0] = t_178[`QUAN_SIZE-1:0];
		`IB_ADDR'd179: t_c[`QUAN_SIZE-1:0] = t_179[`QUAN_SIZE-1:0];
		`IB_ADDR'd180: t_c[`QUAN_SIZE-1:0] = t_180[`QUAN_SIZE-1:0];
		`IB_ADDR'd181: t_c[`QUAN_SIZE-1:0] = t_181[`QUAN_SIZE-1:0];
		`IB_ADDR'd182: t_c[`QUAN_SIZE-1:0] = t_182[`QUAN_SIZE-1:0];
		`IB_ADDR'd183: t_c[`QUAN_SIZE-1:0] = t_183[`QUAN_SIZE-1:0];
		`IB_ADDR'd184: t_c[`QUAN_SIZE-1:0] = t_184[`QUAN_SIZE-1:0];
		`IB_ADDR'd185: t_c[`QUAN_SIZE-1:0] = t_185[`QUAN_SIZE-1:0];
		`IB_ADDR'd186: t_c[`QUAN_SIZE-1:0] = t_186[`QUAN_SIZE-1:0];
		`IB_ADDR'd187: t_c[`QUAN_SIZE-1:0] = t_187[`QUAN_SIZE-1:0];
		`IB_ADDR'd188: t_c[`QUAN_SIZE-1:0] = t_188[`QUAN_SIZE-1:0];
		`IB_ADDR'd189: t_c[`QUAN_SIZE-1:0] = t_189[`QUAN_SIZE-1:0];
		`IB_ADDR'd190: t_c[`QUAN_SIZE-1:0] = t_190[`QUAN_SIZE-1:0];
		`IB_ADDR'd191: t_c[`QUAN_SIZE-1:0] = t_191[`QUAN_SIZE-1:0];
		`IB_ADDR'd192: t_c[`QUAN_SIZE-1:0] = t_192[`QUAN_SIZE-1:0];
		`IB_ADDR'd193: t_c[`QUAN_SIZE-1:0] = t_193[`QUAN_SIZE-1:0];
		`IB_ADDR'd194: t_c[`QUAN_SIZE-1:0] = t_194[`QUAN_SIZE-1:0];
		`IB_ADDR'd195: t_c[`QUAN_SIZE-1:0] = t_195[`QUAN_SIZE-1:0];
		`IB_ADDR'd196: t_c[`QUAN_SIZE-1:0] = t_196[`QUAN_SIZE-1:0];
		`IB_ADDR'd197: t_c[`QUAN_SIZE-1:0] = t_197[`QUAN_SIZE-1:0];
		`IB_ADDR'd198: t_c[`QUAN_SIZE-1:0] = t_198[`QUAN_SIZE-1:0];
		`IB_ADDR'd199: t_c[`QUAN_SIZE-1:0] = t_199[`QUAN_SIZE-1:0];
		`IB_ADDR'd200: t_c[`QUAN_SIZE-1:0] = t_200[`QUAN_SIZE-1:0];
		`IB_ADDR'd201: t_c[`QUAN_SIZE-1:0] = t_201[`QUAN_SIZE-1:0];
		`IB_ADDR'd202: t_c[`QUAN_SIZE-1:0] = t_202[`QUAN_SIZE-1:0];
		`IB_ADDR'd203: t_c[`QUAN_SIZE-1:0] = t_203[`QUAN_SIZE-1:0];
		`IB_ADDR'd204: t_c[`QUAN_SIZE-1:0] = t_204[`QUAN_SIZE-1:0];
		`IB_ADDR'd205: t_c[`QUAN_SIZE-1:0] = t_205[`QUAN_SIZE-1:0];
		`IB_ADDR'd206: t_c[`QUAN_SIZE-1:0] = t_206[`QUAN_SIZE-1:0];
		`IB_ADDR'd207: t_c[`QUAN_SIZE-1:0] = t_207[`QUAN_SIZE-1:0];
		`IB_ADDR'd208: t_c[`QUAN_SIZE-1:0] = t_208[`QUAN_SIZE-1:0];
		`IB_ADDR'd209: t_c[`QUAN_SIZE-1:0] = t_209[`QUAN_SIZE-1:0];
		`IB_ADDR'd210: t_c[`QUAN_SIZE-1:0] = t_210[`QUAN_SIZE-1:0];
		`IB_ADDR'd211: t_c[`QUAN_SIZE-1:0] = t_211[`QUAN_SIZE-1:0];
		`IB_ADDR'd212: t_c[`QUAN_SIZE-1:0] = t_212[`QUAN_SIZE-1:0];
		`IB_ADDR'd213: t_c[`QUAN_SIZE-1:0] = t_213[`QUAN_SIZE-1:0];
		`IB_ADDR'd214: t_c[`QUAN_SIZE-1:0] = t_214[`QUAN_SIZE-1:0];
		`IB_ADDR'd215: t_c[`QUAN_SIZE-1:0] = t_215[`QUAN_SIZE-1:0];
		`IB_ADDR'd216: t_c[`QUAN_SIZE-1:0] = t_216[`QUAN_SIZE-1:0];
		`IB_ADDR'd217: t_c[`QUAN_SIZE-1:0] = t_217[`QUAN_SIZE-1:0];
		`IB_ADDR'd218: t_c[`QUAN_SIZE-1:0] = t_218[`QUAN_SIZE-1:0];
		`IB_ADDR'd219: t_c[`QUAN_SIZE-1:0] = t_219[`QUAN_SIZE-1:0];
		`IB_ADDR'd220: t_c[`QUAN_SIZE-1:0] = t_220[`QUAN_SIZE-1:0];
		`IB_ADDR'd221: t_c[`QUAN_SIZE-1:0] = t_221[`QUAN_SIZE-1:0];
		`IB_ADDR'd222: t_c[`QUAN_SIZE-1:0] = t_222[`QUAN_SIZE-1:0];
		`IB_ADDR'd223: t_c[`QUAN_SIZE-1:0] = t_223[`QUAN_SIZE-1:0];
		`IB_ADDR'd224: t_c[`QUAN_SIZE-1:0] = t_224[`QUAN_SIZE-1:0];
		`IB_ADDR'd225: t_c[`QUAN_SIZE-1:0] = t_225[`QUAN_SIZE-1:0];
		`IB_ADDR'd226: t_c[`QUAN_SIZE-1:0] = t_226[`QUAN_SIZE-1:0];
		`IB_ADDR'd227: t_c[`QUAN_SIZE-1:0] = t_227[`QUAN_SIZE-1:0];
		`IB_ADDR'd228: t_c[`QUAN_SIZE-1:0] = t_228[`QUAN_SIZE-1:0];
		`IB_ADDR'd229: t_c[`QUAN_SIZE-1:0] = t_229[`QUAN_SIZE-1:0];
		`IB_ADDR'd230: t_c[`QUAN_SIZE-1:0] = t_230[`QUAN_SIZE-1:0];
		`IB_ADDR'd231: t_c[`QUAN_SIZE-1:0] = t_231[`QUAN_SIZE-1:0];
		`IB_ADDR'd232: t_c[`QUAN_SIZE-1:0] = t_232[`QUAN_SIZE-1:0];
		`IB_ADDR'd233: t_c[`QUAN_SIZE-1:0] = t_233[`QUAN_SIZE-1:0];
		`IB_ADDR'd234: t_c[`QUAN_SIZE-1:0] = t_234[`QUAN_SIZE-1:0];
		`IB_ADDR'd235: t_c[`QUAN_SIZE-1:0] = t_235[`QUAN_SIZE-1:0];
		`IB_ADDR'd236: t_c[`QUAN_SIZE-1:0] = t_236[`QUAN_SIZE-1:0];
		`IB_ADDR'd237: t_c[`QUAN_SIZE-1:0] = t_237[`QUAN_SIZE-1:0];
		`IB_ADDR'd238: t_c[`QUAN_SIZE-1:0] = t_238[`QUAN_SIZE-1:0];
		`IB_ADDR'd239: t_c[`QUAN_SIZE-1:0] = t_239[`QUAN_SIZE-1:0];
		`IB_ADDR'd240: t_c[`QUAN_SIZE-1:0] = t_240[`QUAN_SIZE-1:0];
		`IB_ADDR'd241: t_c[`QUAN_SIZE-1:0] = t_241[`QUAN_SIZE-1:0];
		`IB_ADDR'd242: t_c[`QUAN_SIZE-1:0] = t_242[`QUAN_SIZE-1:0];
		`IB_ADDR'd243: t_c[`QUAN_SIZE-1:0] = t_243[`QUAN_SIZE-1:0];
		`IB_ADDR'd244: t_c[`QUAN_SIZE-1:0] = t_244[`QUAN_SIZE-1:0];
		`IB_ADDR'd245: t_c[`QUAN_SIZE-1:0] = t_245[`QUAN_SIZE-1:0];
		`IB_ADDR'd246: t_c[`QUAN_SIZE-1:0] = t_246[`QUAN_SIZE-1:0];
		`IB_ADDR'd247: t_c[`QUAN_SIZE-1:0] = t_247[`QUAN_SIZE-1:0];
		`IB_ADDR'd248: t_c[`QUAN_SIZE-1:0] = t_248[`QUAN_SIZE-1:0];
		`IB_ADDR'd249: t_c[`QUAN_SIZE-1:0] = t_249[`QUAN_SIZE-1:0];
		`IB_ADDR'd250: t_c[`QUAN_SIZE-1:0] = t_250[`QUAN_SIZE-1:0];
		`IB_ADDR'd251: t_c[`QUAN_SIZE-1:0] = t_251[`QUAN_SIZE-1:0];
		`IB_ADDR'd252: t_c[`QUAN_SIZE-1:0] = t_252[`QUAN_SIZE-1:0];
		`IB_ADDR'd253: t_c[`QUAN_SIZE-1:0] = t_253[`QUAN_SIZE-1:0];
		`IB_ADDR'd254: t_c[`QUAN_SIZE-1:0] = t_254[`QUAN_SIZE-1:0];
		`IB_ADDR'd255: t_c[`QUAN_SIZE-1:0] = t_255[`QUAN_SIZE-1:0];
	endcase
end
endmodule
