always @(posedge sys_clk) begin
	case(addr_in[`IB_ADDR-1:0])
		`IB_ADDR'd0t_c[`QUAN_SIZE-1:0] <= t_0[`QUAN_SIZE-1:0];
		`IB_ADDR'd1t_c[`QUAN_SIZE-1:0] <= t_1[`QUAN_SIZE-1:0];
		`IB_ADDR'd2t_c[`QUAN_SIZE-1:0] <= t_2[`QUAN_SIZE-1:0];
		`IB_ADDR'd3t_c[`QUAN_SIZE-1:0] <= t_3[`QUAN_SIZE-1:0];
		`IB_ADDR'd4t_c[`QUAN_SIZE-1:0] <= t_4[`QUAN_SIZE-1:0];
		`IB_ADDR'd5t_c[`QUAN_SIZE-1:0] <= t_5[`QUAN_SIZE-1:0];
		`IB_ADDR'd6t_c[`QUAN_SIZE-1:0] <= t_6[`QUAN_SIZE-1:0];
		`IB_ADDR'd7t_c[`QUAN_SIZE-1:0] <= t_7[`QUAN_SIZE-1:0];
		`IB_ADDR'd8t_c[`QUAN_SIZE-1:0] <= t_8[`QUAN_SIZE-1:0];
		`IB_ADDR'd9t_c[`QUAN_SIZE-1:0] <= t_9[`QUAN_SIZE-1:0];
		`IB_ADDR'd10t_c[`QUAN_SIZE-1:0] <= t_10[`QUAN_SIZE-1:0];
		`IB_ADDR'd11t_c[`QUAN_SIZE-1:0] <= t_11[`QUAN_SIZE-1:0];
		`IB_ADDR'd12t_c[`QUAN_SIZE-1:0] <= t_12[`QUAN_SIZE-1:0];
		`IB_ADDR'd13t_c[`QUAN_SIZE-1:0] <= t_13[`QUAN_SIZE-1:0];
		`IB_ADDR'd14t_c[`QUAN_SIZE-1:0] <= t_14[`QUAN_SIZE-1:0];
		`IB_ADDR'd15t_c[`QUAN_SIZE-1:0] <= t_15[`QUAN_SIZE-1:0];
		`IB_ADDR'd16t_c[`QUAN_SIZE-1:0] <= t_16[`QUAN_SIZE-1:0];
		`IB_ADDR'd17t_c[`QUAN_SIZE-1:0] <= t_17[`QUAN_SIZE-1:0];
		`IB_ADDR'd18t_c[`QUAN_SIZE-1:0] <= t_18[`QUAN_SIZE-1:0];
		`IB_ADDR'd19t_c[`QUAN_SIZE-1:0] <= t_19[`QUAN_SIZE-1:0];
		`IB_ADDR'd20t_c[`QUAN_SIZE-1:0] <= t_20[`QUAN_SIZE-1:0];
		`IB_ADDR'd21t_c[`QUAN_SIZE-1:0] <= t_21[`QUAN_SIZE-1:0];
		`IB_ADDR'd22t_c[`QUAN_SIZE-1:0] <= t_22[`QUAN_SIZE-1:0];
		`IB_ADDR'd23t_c[`QUAN_SIZE-1:0] <= t_23[`QUAN_SIZE-1:0];
		`IB_ADDR'd24t_c[`QUAN_SIZE-1:0] <= t_24[`QUAN_SIZE-1:0];
		`IB_ADDR'd25t_c[`QUAN_SIZE-1:0] <= t_25[`QUAN_SIZE-1:0];
		`IB_ADDR'd26t_c[`QUAN_SIZE-1:0] <= t_26[`QUAN_SIZE-1:0];
		`IB_ADDR'd27t_c[`QUAN_SIZE-1:0] <= t_27[`QUAN_SIZE-1:0];
		`IB_ADDR'd28t_c[`QUAN_SIZE-1:0] <= t_28[`QUAN_SIZE-1:0];
		`IB_ADDR'd29t_c[`QUAN_SIZE-1:0] <= t_29[`QUAN_SIZE-1:0];
		`IB_ADDR'd30t_c[`QUAN_SIZE-1:0] <= t_30[`QUAN_SIZE-1:0];
		`IB_ADDR'd31t_c[`QUAN_SIZE-1:0] <= t_31[`QUAN_SIZE-1:0];
		`IB_ADDR'd32t_c[`QUAN_SIZE-1:0] <= t_32[`QUAN_SIZE-1:0];
		`IB_ADDR'd33t_c[`QUAN_SIZE-1:0] <= t_33[`QUAN_SIZE-1:0];
		`IB_ADDR'd34t_c[`QUAN_SIZE-1:0] <= t_34[`QUAN_SIZE-1:0];
		`IB_ADDR'd35t_c[`QUAN_SIZE-1:0] <= t_35[`QUAN_SIZE-1:0];
		`IB_ADDR'd36t_c[`QUAN_SIZE-1:0] <= t_36[`QUAN_SIZE-1:0];
		`IB_ADDR'd37t_c[`QUAN_SIZE-1:0] <= t_37[`QUAN_SIZE-1:0];
		`IB_ADDR'd38t_c[`QUAN_SIZE-1:0] <= t_38[`QUAN_SIZE-1:0];
		`IB_ADDR'd39t_c[`QUAN_SIZE-1:0] <= t_39[`QUAN_SIZE-1:0];
		`IB_ADDR'd40t_c[`QUAN_SIZE-1:0] <= t_40[`QUAN_SIZE-1:0];
		`IB_ADDR'd41t_c[`QUAN_SIZE-1:0] <= t_41[`QUAN_SIZE-1:0];
		`IB_ADDR'd42t_c[`QUAN_SIZE-1:0] <= t_42[`QUAN_SIZE-1:0];
		`IB_ADDR'd43t_c[`QUAN_SIZE-1:0] <= t_43[`QUAN_SIZE-1:0];
		`IB_ADDR'd44t_c[`QUAN_SIZE-1:0] <= t_44[`QUAN_SIZE-1:0];
		`IB_ADDR'd45t_c[`QUAN_SIZE-1:0] <= t_45[`QUAN_SIZE-1:0];
		`IB_ADDR'd46t_c[`QUAN_SIZE-1:0] <= t_46[`QUAN_SIZE-1:0];
		`IB_ADDR'd47t_c[`QUAN_SIZE-1:0] <= t_47[`QUAN_SIZE-1:0];
		`IB_ADDR'd48t_c[`QUAN_SIZE-1:0] <= t_48[`QUAN_SIZE-1:0];
		`IB_ADDR'd49t_c[`QUAN_SIZE-1:0] <= t_49[`QUAN_SIZE-1:0];
		`IB_ADDR'd50t_c[`QUAN_SIZE-1:0] <= t_50[`QUAN_SIZE-1:0];
		`IB_ADDR'd51t_c[`QUAN_SIZE-1:0] <= t_51[`QUAN_SIZE-1:0];
		`IB_ADDR'd52t_c[`QUAN_SIZE-1:0] <= t_52[`QUAN_SIZE-1:0];
		`IB_ADDR'd53t_c[`QUAN_SIZE-1:0] <= t_53[`QUAN_SIZE-1:0];
		`IB_ADDR'd54t_c[`QUAN_SIZE-1:0] <= t_54[`QUAN_SIZE-1:0];
		`IB_ADDR'd55t_c[`QUAN_SIZE-1:0] <= t_55[`QUAN_SIZE-1:0];
		`IB_ADDR'd56t_c[`QUAN_SIZE-1:0] <= t_56[`QUAN_SIZE-1:0];
		`IB_ADDR'd57t_c[`QUAN_SIZE-1:0] <= t_57[`QUAN_SIZE-1:0];
		`IB_ADDR'd58t_c[`QUAN_SIZE-1:0] <= t_58[`QUAN_SIZE-1:0];
		`IB_ADDR'd59t_c[`QUAN_SIZE-1:0] <= t_59[`QUAN_SIZE-1:0];
		`IB_ADDR'd60t_c[`QUAN_SIZE-1:0] <= t_60[`QUAN_SIZE-1:0];
		`IB_ADDR'd61t_c[`QUAN_SIZE-1:0] <= t_61[`QUAN_SIZE-1:0];
		`IB_ADDR'd62t_c[`QUAN_SIZE-1:0] <= t_62[`QUAN_SIZE-1:0];
		`IB_ADDR'd63t_c[`QUAN_SIZE-1:0] <= t_63[`QUAN_SIZE-1:0];
		`IB_ADDR'd64t_c[`QUAN_SIZE-1:0] <= t_64[`QUAN_SIZE-1:0];
		`IB_ADDR'd65t_c[`QUAN_SIZE-1:0] <= t_65[`QUAN_SIZE-1:0];
		`IB_ADDR'd66t_c[`QUAN_SIZE-1:0] <= t_66[`QUAN_SIZE-1:0];
		`IB_ADDR'd67t_c[`QUAN_SIZE-1:0] <= t_67[`QUAN_SIZE-1:0];
		`IB_ADDR'd68t_c[`QUAN_SIZE-1:0] <= t_68[`QUAN_SIZE-1:0];
		`IB_ADDR'd69t_c[`QUAN_SIZE-1:0] <= t_69[`QUAN_SIZE-1:0];
		`IB_ADDR'd70t_c[`QUAN_SIZE-1:0] <= t_70[`QUAN_SIZE-1:0];
		`IB_ADDR'd71t_c[`QUAN_SIZE-1:0] <= t_71[`QUAN_SIZE-1:0];
		`IB_ADDR'd72t_c[`QUAN_SIZE-1:0] <= t_72[`QUAN_SIZE-1:0];
		`IB_ADDR'd73t_c[`QUAN_SIZE-1:0] <= t_73[`QUAN_SIZE-1:0];
		`IB_ADDR'd74t_c[`QUAN_SIZE-1:0] <= t_74[`QUAN_SIZE-1:0];
		`IB_ADDR'd75t_c[`QUAN_SIZE-1:0] <= t_75[`QUAN_SIZE-1:0];
		`IB_ADDR'd76t_c[`QUAN_SIZE-1:0] <= t_76[`QUAN_SIZE-1:0];
		`IB_ADDR'd77t_c[`QUAN_SIZE-1:0] <= t_77[`QUAN_SIZE-1:0];
		`IB_ADDR'd78t_c[`QUAN_SIZE-1:0] <= t_78[`QUAN_SIZE-1:0];
		`IB_ADDR'd79t_c[`QUAN_SIZE-1:0] <= t_79[`QUAN_SIZE-1:0];
		`IB_ADDR'd80t_c[`QUAN_SIZE-1:0] <= t_80[`QUAN_SIZE-1:0];
		`IB_ADDR'd81t_c[`QUAN_SIZE-1:0] <= t_81[`QUAN_SIZE-1:0];
		`IB_ADDR'd82t_c[`QUAN_SIZE-1:0] <= t_82[`QUAN_SIZE-1:0];
		`IB_ADDR'd83t_c[`QUAN_SIZE-1:0] <= t_83[`QUAN_SIZE-1:0];
		`IB_ADDR'd84t_c[`QUAN_SIZE-1:0] <= t_84[`QUAN_SIZE-1:0];
		`IB_ADDR'd85t_c[`QUAN_SIZE-1:0] <= t_85[`QUAN_SIZE-1:0];
		`IB_ADDR'd86t_c[`QUAN_SIZE-1:0] <= t_86[`QUAN_SIZE-1:0];
		`IB_ADDR'd87t_c[`QUAN_SIZE-1:0] <= t_87[`QUAN_SIZE-1:0];
		`IB_ADDR'd88t_c[`QUAN_SIZE-1:0] <= t_88[`QUAN_SIZE-1:0];
		`IB_ADDR'd89t_c[`QUAN_SIZE-1:0] <= t_89[`QUAN_SIZE-1:0];
		`IB_ADDR'd90t_c[`QUAN_SIZE-1:0] <= t_90[`QUAN_SIZE-1:0];
		`IB_ADDR'd91t_c[`QUAN_SIZE-1:0] <= t_91[`QUAN_SIZE-1:0];
		`IB_ADDR'd92t_c[`QUAN_SIZE-1:0] <= t_92[`QUAN_SIZE-1:0];
		`IB_ADDR'd93t_c[`QUAN_SIZE-1:0] <= t_93[`QUAN_SIZE-1:0];
		`IB_ADDR'd94t_c[`QUAN_SIZE-1:0] <= t_94[`QUAN_SIZE-1:0];
		`IB_ADDR'd95t_c[`QUAN_SIZE-1:0] <= t_95[`QUAN_SIZE-1:0];
		`IB_ADDR'd96t_c[`QUAN_SIZE-1:0] <= t_96[`QUAN_SIZE-1:0];
		`IB_ADDR'd97t_c[`QUAN_SIZE-1:0] <= t_97[`QUAN_SIZE-1:0];
		`IB_ADDR'd98t_c[`QUAN_SIZE-1:0] <= t_98[`QUAN_SIZE-1:0];
		`IB_ADDR'd99t_c[`QUAN_SIZE-1:0] <= t_99[`QUAN_SIZE-1:0];
		`IB_ADDR'd100t_c[`QUAN_SIZE-1:0] <= t_100[`QUAN_SIZE-1:0];
		`IB_ADDR'd101t_c[`QUAN_SIZE-1:0] <= t_101[`QUAN_SIZE-1:0];
		`IB_ADDR'd102t_c[`QUAN_SIZE-1:0] <= t_102[`QUAN_SIZE-1:0];
		`IB_ADDR'd103t_c[`QUAN_SIZE-1:0] <= t_103[`QUAN_SIZE-1:0];
		`IB_ADDR'd104t_c[`QUAN_SIZE-1:0] <= t_104[`QUAN_SIZE-1:0];
		`IB_ADDR'd105t_c[`QUAN_SIZE-1:0] <= t_105[`QUAN_SIZE-1:0];
		`IB_ADDR'd106t_c[`QUAN_SIZE-1:0] <= t_106[`QUAN_SIZE-1:0];
		`IB_ADDR'd107t_c[`QUAN_SIZE-1:0] <= t_107[`QUAN_SIZE-1:0];
		`IB_ADDR'd108t_c[`QUAN_SIZE-1:0] <= t_108[`QUAN_SIZE-1:0];
		`IB_ADDR'd109t_c[`QUAN_SIZE-1:0] <= t_109[`QUAN_SIZE-1:0];
		`IB_ADDR'd110t_c[`QUAN_SIZE-1:0] <= t_110[`QUAN_SIZE-1:0];
		`IB_ADDR'd111t_c[`QUAN_SIZE-1:0] <= t_111[`QUAN_SIZE-1:0];
		`IB_ADDR'd112t_c[`QUAN_SIZE-1:0] <= t_112[`QUAN_SIZE-1:0];
		`IB_ADDR'd113t_c[`QUAN_SIZE-1:0] <= t_113[`QUAN_SIZE-1:0];
		`IB_ADDR'd114t_c[`QUAN_SIZE-1:0] <= t_114[`QUAN_SIZE-1:0];
		`IB_ADDR'd115t_c[`QUAN_SIZE-1:0] <= t_115[`QUAN_SIZE-1:0];
		`IB_ADDR'd116t_c[`QUAN_SIZE-1:0] <= t_116[`QUAN_SIZE-1:0];
		`IB_ADDR'd117t_c[`QUAN_SIZE-1:0] <= t_117[`QUAN_SIZE-1:0];
		`IB_ADDR'd118t_c[`QUAN_SIZE-1:0] <= t_118[`QUAN_SIZE-1:0];
		`IB_ADDR'd119t_c[`QUAN_SIZE-1:0] <= t_119[`QUAN_SIZE-1:0];
		`IB_ADDR'd120t_c[`QUAN_SIZE-1:0] <= t_120[`QUAN_SIZE-1:0];
		`IB_ADDR'd121t_c[`QUAN_SIZE-1:0] <= t_121[`QUAN_SIZE-1:0];
		`IB_ADDR'd122t_c[`QUAN_SIZE-1:0] <= t_122[`QUAN_SIZE-1:0];
		`IB_ADDR'd123t_c[`QUAN_SIZE-1:0] <= t_123[`QUAN_SIZE-1:0];
		`IB_ADDR'd124t_c[`QUAN_SIZE-1:0] <= t_124[`QUAN_SIZE-1:0];
		`IB_ADDR'd125t_c[`QUAN_SIZE-1:0] <= t_125[`QUAN_SIZE-1:0];
		`IB_ADDR'd126t_c[`QUAN_SIZE-1:0] <= t_126[`QUAN_SIZE-1:0];
		`IB_ADDR'd127t_c[`QUAN_SIZE-1:0] <= t_127[`QUAN_SIZE-1:0];
		`IB_ADDR'd128t_c[`QUAN_SIZE-1:0] <= t_128[`QUAN_SIZE-1:0];
		`IB_ADDR'd129t_c[`QUAN_SIZE-1:0] <= t_129[`QUAN_SIZE-1:0];
		`IB_ADDR'd130t_c[`QUAN_SIZE-1:0] <= t_130[`QUAN_SIZE-1:0];
		`IB_ADDR'd131t_c[`QUAN_SIZE-1:0] <= t_131[`QUAN_SIZE-1:0];
		`IB_ADDR'd132t_c[`QUAN_SIZE-1:0] <= t_132[`QUAN_SIZE-1:0];
		`IB_ADDR'd133t_c[`QUAN_SIZE-1:0] <= t_133[`QUAN_SIZE-1:0];
		`IB_ADDR'd134t_c[`QUAN_SIZE-1:0] <= t_134[`QUAN_SIZE-1:0];
		`IB_ADDR'd135t_c[`QUAN_SIZE-1:0] <= t_135[`QUAN_SIZE-1:0];
		`IB_ADDR'd136t_c[`QUAN_SIZE-1:0] <= t_136[`QUAN_SIZE-1:0];
		`IB_ADDR'd137t_c[`QUAN_SIZE-1:0] <= t_137[`QUAN_SIZE-1:0];
		`IB_ADDR'd138t_c[`QUAN_SIZE-1:0] <= t_138[`QUAN_SIZE-1:0];
		`IB_ADDR'd139t_c[`QUAN_SIZE-1:0] <= t_139[`QUAN_SIZE-1:0];
		`IB_ADDR'd140t_c[`QUAN_SIZE-1:0] <= t_140[`QUAN_SIZE-1:0];
		`IB_ADDR'd141t_c[`QUAN_SIZE-1:0] <= t_141[`QUAN_SIZE-1:0];
		`IB_ADDR'd142t_c[`QUAN_SIZE-1:0] <= t_142[`QUAN_SIZE-1:0];
		`IB_ADDR'd143t_c[`QUAN_SIZE-1:0] <= t_143[`QUAN_SIZE-1:0];
		`IB_ADDR'd144t_c[`QUAN_SIZE-1:0] <= t_144[`QUAN_SIZE-1:0];
		`IB_ADDR'd145t_c[`QUAN_SIZE-1:0] <= t_145[`QUAN_SIZE-1:0];
		`IB_ADDR'd146t_c[`QUAN_SIZE-1:0] <= t_146[`QUAN_SIZE-1:0];
		`IB_ADDR'd147t_c[`QUAN_SIZE-1:0] <= t_147[`QUAN_SIZE-1:0];
		`IB_ADDR'd148t_c[`QUAN_SIZE-1:0] <= t_148[`QUAN_SIZE-1:0];
		`IB_ADDR'd149t_c[`QUAN_SIZE-1:0] <= t_149[`QUAN_SIZE-1:0];
		`IB_ADDR'd150t_c[`QUAN_SIZE-1:0] <= t_150[`QUAN_SIZE-1:0];
		`IB_ADDR'd151t_c[`QUAN_SIZE-1:0] <= t_151[`QUAN_SIZE-1:0];
		`IB_ADDR'd152t_c[`QUAN_SIZE-1:0] <= t_152[`QUAN_SIZE-1:0];
		`IB_ADDR'd153t_c[`QUAN_SIZE-1:0] <= t_153[`QUAN_SIZE-1:0];
		`IB_ADDR'd154t_c[`QUAN_SIZE-1:0] <= t_154[`QUAN_SIZE-1:0];
		`IB_ADDR'd155t_c[`QUAN_SIZE-1:0] <= t_155[`QUAN_SIZE-1:0];
		`IB_ADDR'd156t_c[`QUAN_SIZE-1:0] <= t_156[`QUAN_SIZE-1:0];
		`IB_ADDR'd157t_c[`QUAN_SIZE-1:0] <= t_157[`QUAN_SIZE-1:0];
		`IB_ADDR'd158t_c[`QUAN_SIZE-1:0] <= t_158[`QUAN_SIZE-1:0];
		`IB_ADDR'd159t_c[`QUAN_SIZE-1:0] <= t_159[`QUAN_SIZE-1:0];
		`IB_ADDR'd160t_c[`QUAN_SIZE-1:0] <= t_160[`QUAN_SIZE-1:0];
		`IB_ADDR'd161t_c[`QUAN_SIZE-1:0] <= t_161[`QUAN_SIZE-1:0];
		`IB_ADDR'd162t_c[`QUAN_SIZE-1:0] <= t_162[`QUAN_SIZE-1:0];
		`IB_ADDR'd163t_c[`QUAN_SIZE-1:0] <= t_163[`QUAN_SIZE-1:0];
		`IB_ADDR'd164t_c[`QUAN_SIZE-1:0] <= t_164[`QUAN_SIZE-1:0];
		`IB_ADDR'd165t_c[`QUAN_SIZE-1:0] <= t_165[`QUAN_SIZE-1:0];
		`IB_ADDR'd166t_c[`QUAN_SIZE-1:0] <= t_166[`QUAN_SIZE-1:0];
		`IB_ADDR'd167t_c[`QUAN_SIZE-1:0] <= t_167[`QUAN_SIZE-1:0];
		`IB_ADDR'd168t_c[`QUAN_SIZE-1:0] <= t_168[`QUAN_SIZE-1:0];
		`IB_ADDR'd169t_c[`QUAN_SIZE-1:0] <= t_169[`QUAN_SIZE-1:0];
		`IB_ADDR'd170t_c[`QUAN_SIZE-1:0] <= t_170[`QUAN_SIZE-1:0];
		`IB_ADDR'd171t_c[`QUAN_SIZE-1:0] <= t_171[`QUAN_SIZE-1:0];
		`IB_ADDR'd172t_c[`QUAN_SIZE-1:0] <= t_172[`QUAN_SIZE-1:0];
		`IB_ADDR'd173t_c[`QUAN_SIZE-1:0] <= t_173[`QUAN_SIZE-1:0];
		`IB_ADDR'd174t_c[`QUAN_SIZE-1:0] <= t_174[`QUAN_SIZE-1:0];
		`IB_ADDR'd175t_c[`QUAN_SIZE-1:0] <= t_175[`QUAN_SIZE-1:0];
		`IB_ADDR'd176t_c[`QUAN_SIZE-1:0] <= t_176[`QUAN_SIZE-1:0];
		`IB_ADDR'd177t_c[`QUAN_SIZE-1:0] <= t_177[`QUAN_SIZE-1:0];
		`IB_ADDR'd178t_c[`QUAN_SIZE-1:0] <= t_178[`QUAN_SIZE-1:0];
		`IB_ADDR'd179t_c[`QUAN_SIZE-1:0] <= t_179[`QUAN_SIZE-1:0];
		`IB_ADDR'd180t_c[`QUAN_SIZE-1:0] <= t_180[`QUAN_SIZE-1:0];
		`IB_ADDR'd181t_c[`QUAN_SIZE-1:0] <= t_181[`QUAN_SIZE-1:0];
		`IB_ADDR'd182t_c[`QUAN_SIZE-1:0] <= t_182[`QUAN_SIZE-1:0];
		`IB_ADDR'd183t_c[`QUAN_SIZE-1:0] <= t_183[`QUAN_SIZE-1:0];
		`IB_ADDR'd184t_c[`QUAN_SIZE-1:0] <= t_184[`QUAN_SIZE-1:0];
		`IB_ADDR'd185t_c[`QUAN_SIZE-1:0] <= t_185[`QUAN_SIZE-1:0];
		`IB_ADDR'd186t_c[`QUAN_SIZE-1:0] <= t_186[`QUAN_SIZE-1:0];
		`IB_ADDR'd187t_c[`QUAN_SIZE-1:0] <= t_187[`QUAN_SIZE-1:0];
		`IB_ADDR'd188t_c[`QUAN_SIZE-1:0] <= t_188[`QUAN_SIZE-1:0];
		`IB_ADDR'd189t_c[`QUAN_SIZE-1:0] <= t_189[`QUAN_SIZE-1:0];
		`IB_ADDR'd190t_c[`QUAN_SIZE-1:0] <= t_190[`QUAN_SIZE-1:0];
		`IB_ADDR'd191t_c[`QUAN_SIZE-1:0] <= t_191[`QUAN_SIZE-1:0];
		`IB_ADDR'd192t_c[`QUAN_SIZE-1:0] <= t_192[`QUAN_SIZE-1:0];
		`IB_ADDR'd193t_c[`QUAN_SIZE-1:0] <= t_193[`QUAN_SIZE-1:0];
		`IB_ADDR'd194t_c[`QUAN_SIZE-1:0] <= t_194[`QUAN_SIZE-1:0];
		`IB_ADDR'd195t_c[`QUAN_SIZE-1:0] <= t_195[`QUAN_SIZE-1:0];
		`IB_ADDR'd196t_c[`QUAN_SIZE-1:0] <= t_196[`QUAN_SIZE-1:0];
		`IB_ADDR'd197t_c[`QUAN_SIZE-1:0] <= t_197[`QUAN_SIZE-1:0];
		`IB_ADDR'd198t_c[`QUAN_SIZE-1:0] <= t_198[`QUAN_SIZE-1:0];
		`IB_ADDR'd199t_c[`QUAN_SIZE-1:0] <= t_199[`QUAN_SIZE-1:0];
		`IB_ADDR'd200t_c[`QUAN_SIZE-1:0] <= t_200[`QUAN_SIZE-1:0];
		`IB_ADDR'd201t_c[`QUAN_SIZE-1:0] <= t_201[`QUAN_SIZE-1:0];
		`IB_ADDR'd202t_c[`QUAN_SIZE-1:0] <= t_202[`QUAN_SIZE-1:0];
		`IB_ADDR'd203t_c[`QUAN_SIZE-1:0] <= t_203[`QUAN_SIZE-1:0];
		`IB_ADDR'd204t_c[`QUAN_SIZE-1:0] <= t_204[`QUAN_SIZE-1:0];
		`IB_ADDR'd205t_c[`QUAN_SIZE-1:0] <= t_205[`QUAN_SIZE-1:0];
		`IB_ADDR'd206t_c[`QUAN_SIZE-1:0] <= t_206[`QUAN_SIZE-1:0];
		`IB_ADDR'd207t_c[`QUAN_SIZE-1:0] <= t_207[`QUAN_SIZE-1:0];
		`IB_ADDR'd208t_c[`QUAN_SIZE-1:0] <= t_208[`QUAN_SIZE-1:0];
		`IB_ADDR'd209t_c[`QUAN_SIZE-1:0] <= t_209[`QUAN_SIZE-1:0];
		`IB_ADDR'd210t_c[`QUAN_SIZE-1:0] <= t_210[`QUAN_SIZE-1:0];
		`IB_ADDR'd211t_c[`QUAN_SIZE-1:0] <= t_211[`QUAN_SIZE-1:0];
		`IB_ADDR'd212t_c[`QUAN_SIZE-1:0] <= t_212[`QUAN_SIZE-1:0];
		`IB_ADDR'd213t_c[`QUAN_SIZE-1:0] <= t_213[`QUAN_SIZE-1:0];
		`IB_ADDR'd214t_c[`QUAN_SIZE-1:0] <= t_214[`QUAN_SIZE-1:0];
		`IB_ADDR'd215t_c[`QUAN_SIZE-1:0] <= t_215[`QUAN_SIZE-1:0];
		`IB_ADDR'd216t_c[`QUAN_SIZE-1:0] <= t_216[`QUAN_SIZE-1:0];
		`IB_ADDR'd217t_c[`QUAN_SIZE-1:0] <= t_217[`QUAN_SIZE-1:0];
		`IB_ADDR'd218t_c[`QUAN_SIZE-1:0] <= t_218[`QUAN_SIZE-1:0];
		`IB_ADDR'd219t_c[`QUAN_SIZE-1:0] <= t_219[`QUAN_SIZE-1:0];
		`IB_ADDR'd220t_c[`QUAN_SIZE-1:0] <= t_220[`QUAN_SIZE-1:0];
		`IB_ADDR'd221t_c[`QUAN_SIZE-1:0] <= t_221[`QUAN_SIZE-1:0];
		`IB_ADDR'd222t_c[`QUAN_SIZE-1:0] <= t_222[`QUAN_SIZE-1:0];
		`IB_ADDR'd223t_c[`QUAN_SIZE-1:0] <= t_223[`QUAN_SIZE-1:0];
		`IB_ADDR'd224t_c[`QUAN_SIZE-1:0] <= t_224[`QUAN_SIZE-1:0];
		`IB_ADDR'd225t_c[`QUAN_SIZE-1:0] <= t_225[`QUAN_SIZE-1:0];
		`IB_ADDR'd226t_c[`QUAN_SIZE-1:0] <= t_226[`QUAN_SIZE-1:0];
		`IB_ADDR'd227t_c[`QUAN_SIZE-1:0] <= t_227[`QUAN_SIZE-1:0];
		`IB_ADDR'd228t_c[`QUAN_SIZE-1:0] <= t_228[`QUAN_SIZE-1:0];
		`IB_ADDR'd229t_c[`QUAN_SIZE-1:0] <= t_229[`QUAN_SIZE-1:0];
		`IB_ADDR'd230t_c[`QUAN_SIZE-1:0] <= t_230[`QUAN_SIZE-1:0];
		`IB_ADDR'd231t_c[`QUAN_SIZE-1:0] <= t_231[`QUAN_SIZE-1:0];
		`IB_ADDR'd232t_c[`QUAN_SIZE-1:0] <= t_232[`QUAN_SIZE-1:0];
		`IB_ADDR'd233t_c[`QUAN_SIZE-1:0] <= t_233[`QUAN_SIZE-1:0];
		`IB_ADDR'd234t_c[`QUAN_SIZE-1:0] <= t_234[`QUAN_SIZE-1:0];
		`IB_ADDR'd235t_c[`QUAN_SIZE-1:0] <= t_235[`QUAN_SIZE-1:0];
		`IB_ADDR'd236t_c[`QUAN_SIZE-1:0] <= t_236[`QUAN_SIZE-1:0];
		`IB_ADDR'd237t_c[`QUAN_SIZE-1:0] <= t_237[`QUAN_SIZE-1:0];
		`IB_ADDR'd238t_c[`QUAN_SIZE-1:0] <= t_238[`QUAN_SIZE-1:0];
		`IB_ADDR'd239t_c[`QUAN_SIZE-1:0] <= t_239[`QUAN_SIZE-1:0];
		`IB_ADDR'd240t_c[`QUAN_SIZE-1:0] <= t_240[`QUAN_SIZE-1:0];
		`IB_ADDR'd241t_c[`QUAN_SIZE-1:0] <= t_241[`QUAN_SIZE-1:0];
		`IB_ADDR'd242t_c[`QUAN_SIZE-1:0] <= t_242[`QUAN_SIZE-1:0];
		`IB_ADDR'd243t_c[`QUAN_SIZE-1:0] <= t_243[`QUAN_SIZE-1:0];
		`IB_ADDR'd244t_c[`QUAN_SIZE-1:0] <= t_244[`QUAN_SIZE-1:0];
		`IB_ADDR'd245t_c[`QUAN_SIZE-1:0] <= t_245[`QUAN_SIZE-1:0];
		`IB_ADDR'd246t_c[`QUAN_SIZE-1:0] <= t_246[`QUAN_SIZE-1:0];
		`IB_ADDR'd247t_c[`QUAN_SIZE-1:0] <= t_247[`QUAN_SIZE-1:0];
		`IB_ADDR'd248t_c[`QUAN_SIZE-1:0] <= t_248[`QUAN_SIZE-1:0];
		`IB_ADDR'd249t_c[`QUAN_SIZE-1:0] <= t_249[`QUAN_SIZE-1:0];
		`IB_ADDR'd250t_c[`QUAN_SIZE-1:0] <= t_250[`QUAN_SIZE-1:0];
		`IB_ADDR'd251t_c[`QUAN_SIZE-1:0] <= t_251[`QUAN_SIZE-1:0];
		`IB_ADDR'd252t_c[`QUAN_SIZE-1:0] <= t_252[`QUAN_SIZE-1:0];
		`IB_ADDR'd253t_c[`QUAN_SIZE-1:0] <= t_253[`QUAN_SIZE-1:0];
		`IB_ADDR'd254t_c[`QUAN_SIZE-1:0] <= t_254[`QUAN_SIZE-1:0];
		`IB_ADDR'd255t_c[`QUAN_SIZE-1:0] <= t_255[`QUAN_SIZE-1:0];
	endcase
end