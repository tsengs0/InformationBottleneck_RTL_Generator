
`timescale 1ns/1ps

module tb_mem_subsystem_top (); /* this is automatically generated */

	// clock
	logic clk;
	initial begin
		clk = '0;
		forever #(0.5) clk = ~clk;
	end

	// synchronous reset
	logic srstb;
	initial begin
		srstb <= '0;
		repeat(10)@(posedge clk);
		srstb <= '1;
	end

	// (*NOTE*) replace reset, clock, others

	parameter         QUAN_SIZE = 4;
	parameter CHECK_PARALLELISM = 85;
	parameter         LAYER_NUM = 3;
	parameter  RAM_UNIT_MSG_NUM = 17;
	parameter   RAM_PORTA_RANGE = 9;
	parameter   RAM_PORTB_RANGE = 8;
	parameter    MEM_DEVICE_NUM = 5;
	parameter             DEPTH = 1024;
	parameter             WIDTH = 36;
	parameter              ADDR = $clog2(DEPTH);

	logic         [QUAN_SIZE-1:0] mem_to_bs_0;
	logic         [QUAN_SIZE-1:0] mem_to_bs_1;
	logic         [QUAN_SIZE-1:0] mem_to_bs_2;
	logic         [QUAN_SIZE-1:0] mem_to_bs_3;
	logic         [QUAN_SIZE-1:0] mem_to_bs_4;
	logic         [QUAN_SIZE-1:0] mem_to_bs_5;
	logic         [QUAN_SIZE-1:0] mem_to_bs_6;
	logic         [QUAN_SIZE-1:0] mem_to_bs_7;
	logic         [QUAN_SIZE-1:0] mem_to_bs_8;
	logic         [QUAN_SIZE-1:0] mem_to_bs_9;
	logic         [QUAN_SIZE-1:0] mem_to_bs_10;
	logic         [QUAN_SIZE-1:0] mem_to_bs_11;
	logic         [QUAN_SIZE-1:0] mem_to_bs_12;
	logic         [QUAN_SIZE-1:0] mem_to_bs_13;
	logic         [QUAN_SIZE-1:0] mem_to_bs_14;
	logic         [QUAN_SIZE-1:0] mem_to_bs_15;
	logic         [QUAN_SIZE-1:0] mem_to_bs_16;
	logic         [QUAN_SIZE-1:0] mem_to_bs_17;
	logic         [QUAN_SIZE-1:0] mem_to_bs_18;
	logic         [QUAN_SIZE-1:0] mem_to_bs_19;
	logic         [QUAN_SIZE-1:0] mem_to_bs_20;
	logic         [QUAN_SIZE-1:0] mem_to_bs_21;
	logic         [QUAN_SIZE-1:0] mem_to_bs_22;
	logic         [QUAN_SIZE-1:0] mem_to_bs_23;
	logic         [QUAN_SIZE-1:0] mem_to_bs_24;
	logic         [QUAN_SIZE-1:0] mem_to_bs_25;
	logic         [QUAN_SIZE-1:0] mem_to_bs_26;
	logic         [QUAN_SIZE-1:0] mem_to_bs_27;
	logic         [QUAN_SIZE-1:0] mem_to_bs_28;
	logic         [QUAN_SIZE-1:0] mem_to_bs_29;
	logic         [QUAN_SIZE-1:0] mem_to_bs_30;
	logic         [QUAN_SIZE-1:0] mem_to_bs_31;
	logic         [QUAN_SIZE-1:0] mem_to_bs_32;
	logic         [QUAN_SIZE-1:0] mem_to_bs_33;
	logic         [QUAN_SIZE-1:0] mem_to_bs_34;
	logic         [QUAN_SIZE-1:0] mem_to_bs_35;
	logic         [QUAN_SIZE-1:0] mem_to_bs_36;
	logic         [QUAN_SIZE-1:0] mem_to_bs_37;
	logic         [QUAN_SIZE-1:0] mem_to_bs_38;
	logic         [QUAN_SIZE-1:0] mem_to_bs_39;
	logic         [QUAN_SIZE-1:0] mem_to_bs_40;
	logic         [QUAN_SIZE-1:0] mem_to_bs_41;
	logic         [QUAN_SIZE-1:0] mem_to_bs_42;
	logic         [QUAN_SIZE-1:0] mem_to_bs_43;
	logic         [QUAN_SIZE-1:0] mem_to_bs_44;
	logic         [QUAN_SIZE-1:0] mem_to_bs_45;
	logic         [QUAN_SIZE-1:0] mem_to_bs_46;
	logic         [QUAN_SIZE-1:0] mem_to_bs_47;
	logic         [QUAN_SIZE-1:0] mem_to_bs_48;
	logic         [QUAN_SIZE-1:0] mem_to_bs_49;
	logic         [QUAN_SIZE-1:0] mem_to_bs_50;
	logic         [QUAN_SIZE-1:0] mem_to_bs_51;
	logic         [QUAN_SIZE-1:0] mem_to_bs_52;
	logic         [QUAN_SIZE-1:0] mem_to_bs_53;
	logic         [QUAN_SIZE-1:0] mem_to_bs_54;
	logic         [QUAN_SIZE-1:0] mem_to_bs_55;
	logic         [QUAN_SIZE-1:0] mem_to_bs_56;
	logic         [QUAN_SIZE-1:0] mem_to_bs_57;
	logic         [QUAN_SIZE-1:0] mem_to_bs_58;
	logic         [QUAN_SIZE-1:0] mem_to_bs_59;
	logic         [QUAN_SIZE-1:0] mem_to_bs_60;
	logic         [QUAN_SIZE-1:0] mem_to_bs_61;
	logic         [QUAN_SIZE-1:0] mem_to_bs_62;
	logic         [QUAN_SIZE-1:0] mem_to_bs_63;
	logic         [QUAN_SIZE-1:0] mem_to_bs_64;
	logic         [QUAN_SIZE-1:0] mem_to_bs_65;
	logic         [QUAN_SIZE-1:0] mem_to_bs_66;
	logic         [QUAN_SIZE-1:0] mem_to_bs_67;
	logic         [QUAN_SIZE-1:0] mem_to_bs_68;
	logic         [QUAN_SIZE-1:0] mem_to_bs_69;
	logic         [QUAN_SIZE-1:0] mem_to_bs_70;
	logic         [QUAN_SIZE-1:0] mem_to_bs_71;
	logic         [QUAN_SIZE-1:0] mem_to_bs_72;
	logic         [QUAN_SIZE-1:0] mem_to_bs_73;
	logic         [QUAN_SIZE-1:0] mem_to_bs_74;
	logic         [QUAN_SIZE-1:0] mem_to_bs_75;
	logic         [QUAN_SIZE-1:0] mem_to_bs_76;
	logic         [QUAN_SIZE-1:0] mem_to_bs_77;
	logic         [QUAN_SIZE-1:0] mem_to_bs_78;
	logic         [QUAN_SIZE-1:0] mem_to_bs_79;
	logic         [QUAN_SIZE-1:0] mem_to_bs_80;
	logic         [QUAN_SIZE-1:0] mem_to_bs_81;
	logic         [QUAN_SIZE-1:0] mem_to_bs_82;
	logic         [QUAN_SIZE-1:0] mem_to_bs_83;
	logic         [QUAN_SIZE-1:0] mem_to_bs_84;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_0;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_1;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_2;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_3;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_4;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_5;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_6;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_7;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_8;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_9;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_10;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_11;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_12;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_13;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_14;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_15;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_16;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_17;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_18;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_19;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_20;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_21;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_22;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_23;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_24;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_25;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_26;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_27;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_28;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_29;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_30;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_31;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_32;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_33;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_34;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_35;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_36;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_37;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_38;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_39;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_40;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_41;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_42;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_43;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_44;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_45;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_46;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_47;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_48;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_49;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_50;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_51;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_52;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_53;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_54;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_55;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_56;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_57;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_58;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_59;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_60;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_61;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_62;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_63;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_64;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_65;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_66;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_67;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_68;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_69;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_70;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_71;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_72;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_73;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_74;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_75;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_76;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_77;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_78;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_79;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_80;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_81;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_82;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_83;
	logic         [QUAN_SIZE-1:0] mem_to_cnu_84;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_1;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_1;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_2;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_3;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_4;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_5;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_6;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_7;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_8;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_9;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_10;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_11;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_12;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_13;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_14;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_15;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_16;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_17;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_18;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_19;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_20;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_21;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_22;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_23;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_24;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_25;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_26;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_27;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_28;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_29;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_30;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_31;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_32;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_33;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_34;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_35;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_36;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_37;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_38;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_39;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_40;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_41;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_42;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_43;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_44;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_45;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_46;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_47;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_48;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_49;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_50;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_51;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_52;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_53;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_54;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_55;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_56;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_57;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_58;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_59;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_60;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_61;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_62;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_63;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_64;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_65;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_66;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_67;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_68;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_69;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_70;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_71;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_72;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_73;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_74;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_75;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_76;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_77;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_78;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_79;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_80;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_81;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_82;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_83;
	logic         [QUAN_SIZE-1:0] vnu_to_mem_84;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_0;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_1;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_2;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_3;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_4;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_5;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_6;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_7;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_8;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_9;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_10;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_11;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_12;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_13;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_14;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_15;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_16;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_17;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_18;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_19;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_20;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_21;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_22;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_23;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_24;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_25;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_26;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_27;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_28;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_29;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_30;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_31;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_32;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_33;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_34;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_35;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_36;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_37;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_38;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_39;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_40;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_41;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_42;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_43;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_44;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_45;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_46;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_47;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_48;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_49;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_50;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_51;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_52;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_53;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_54;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_55;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_56;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_57;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_58;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_59;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_60;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_61;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_62;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_63;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_64;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_65;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_66;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_67;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_68;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_69;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_70;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_71;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_72;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_73;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_74;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_75;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_76;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_77;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_78;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_79;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_80;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_81;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_82;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_83;
	logic         [QUAN_SIZE-1:0] cnu_to_mem_84;
	logic                         sched_cmd;
	logic [CHECK_PARALLELISM-1:0] delay_cmd;
	logic              [ADDR-1:0] sync_addr;
	logic         [LAYER_NUM-1:0] layer_status;
	logic                         first_row_chunk;
	logic                         we;
	logic                         sys_clk;
	logic                         rstn;

	mem_subsystem_top #(
			.QUAN_SIZE(QUAN_SIZE),
			.CHECK_PARALLELISM(CHECK_PARALLELISM),
			.LAYER_NUM(LAYER_NUM),
			.RAM_UNIT_MSG_NUM(RAM_UNIT_MSG_NUM),
			.RAM_PORTA_RANGE(RAM_PORTA_RANGE),
			.RAM_PORTB_RANGE(RAM_PORTB_RANGE),
			.MEM_DEVICE_NUM(MEM_DEVICE_NUM),
			.DEPTH(DEPTH),
			.WIDTH(WIDTH),
			.ADDR(ADDR)
		) inst_mem_subsystem_top (
			.mem_to_bs_0     (mem_to_bs_0),
			.mem_to_bs_1     (mem_to_bs_1),
			.mem_to_bs_2     (mem_to_bs_2),
			.mem_to_bs_3     (mem_to_bs_3),
			.mem_to_bs_4     (mem_to_bs_4),
			.mem_to_bs_5     (mem_to_bs_5),
			.mem_to_bs_6     (mem_to_bs_6),
			.mem_to_bs_7     (mem_to_bs_7),
			.mem_to_bs_8     (mem_to_bs_8),
			.mem_to_bs_9     (mem_to_bs_9),
			.mem_to_bs_10    (mem_to_bs_10),
			.mem_to_bs_11    (mem_to_bs_11),
			.mem_to_bs_12    (mem_to_bs_12),
			.mem_to_bs_13    (mem_to_bs_13),
			.mem_to_bs_14    (mem_to_bs_14),
			.mem_to_bs_15    (mem_to_bs_15),
			.mem_to_bs_16    (mem_to_bs_16),
			.mem_to_bs_17    (mem_to_bs_17),
			.mem_to_bs_18    (mem_to_bs_18),
			.mem_to_bs_19    (mem_to_bs_19),
			.mem_to_bs_20    (mem_to_bs_20),
			.mem_to_bs_21    (mem_to_bs_21),
			.mem_to_bs_22    (mem_to_bs_22),
			.mem_to_bs_23    (mem_to_bs_23),
			.mem_to_bs_24    (mem_to_bs_24),
			.mem_to_bs_25    (mem_to_bs_25),
			.mem_to_bs_26    (mem_to_bs_26),
			.mem_to_bs_27    (mem_to_bs_27),
			.mem_to_bs_28    (mem_to_bs_28),
			.mem_to_bs_29    (mem_to_bs_29),
			.mem_to_bs_30    (mem_to_bs_30),
			.mem_to_bs_31    (mem_to_bs_31),
			.mem_to_bs_32    (mem_to_bs_32),
			.mem_to_bs_33    (mem_to_bs_33),
			.mem_to_bs_34    (mem_to_bs_34),
			.mem_to_bs_35    (mem_to_bs_35),
			.mem_to_bs_36    (mem_to_bs_36),
			.mem_to_bs_37    (mem_to_bs_37),
			.mem_to_bs_38    (mem_to_bs_38),
			.mem_to_bs_39    (mem_to_bs_39),
			.mem_to_bs_40    (mem_to_bs_40),
			.mem_to_bs_41    (mem_to_bs_41),
			.mem_to_bs_42    (mem_to_bs_42),
			.mem_to_bs_43    (mem_to_bs_43),
			.mem_to_bs_44    (mem_to_bs_44),
			.mem_to_bs_45    (mem_to_bs_45),
			.mem_to_bs_46    (mem_to_bs_46),
			.mem_to_bs_47    (mem_to_bs_47),
			.mem_to_bs_48    (mem_to_bs_48),
			.mem_to_bs_49    (mem_to_bs_49),
			.mem_to_bs_50    (mem_to_bs_50),
			.mem_to_bs_51    (mem_to_bs_51),
			.mem_to_bs_52    (mem_to_bs_52),
			.mem_to_bs_53    (mem_to_bs_53),
			.mem_to_bs_54    (mem_to_bs_54),
			.mem_to_bs_55    (mem_to_bs_55),
			.mem_to_bs_56    (mem_to_bs_56),
			.mem_to_bs_57    (mem_to_bs_57),
			.mem_to_bs_58    (mem_to_bs_58),
			.mem_to_bs_59    (mem_to_bs_59),
			.mem_to_bs_60    (mem_to_bs_60),
			.mem_to_bs_61    (mem_to_bs_61),
			.mem_to_bs_62    (mem_to_bs_62),
			.mem_to_bs_63    (mem_to_bs_63),
			.mem_to_bs_64    (mem_to_bs_64),
			.mem_to_bs_65    (mem_to_bs_65),
			.mem_to_bs_66    (mem_to_bs_66),
			.mem_to_bs_67    (mem_to_bs_67),
			.mem_to_bs_68    (mem_to_bs_68),
			.mem_to_bs_69    (mem_to_bs_69),
			.mem_to_bs_70    (mem_to_bs_70),
			.mem_to_bs_71    (mem_to_bs_71),
			.mem_to_bs_72    (mem_to_bs_72),
			.mem_to_bs_73    (mem_to_bs_73),
			.mem_to_bs_74    (mem_to_bs_74),
			.mem_to_bs_75    (mem_to_bs_75),
			.mem_to_bs_76    (mem_to_bs_76),
			.mem_to_bs_77    (mem_to_bs_77),
			.mem_to_bs_78    (mem_to_bs_78),
			.mem_to_bs_79    (mem_to_bs_79),
			.mem_to_bs_80    (mem_to_bs_80),
			.mem_to_bs_81    (mem_to_bs_81),
			.mem_to_bs_82    (mem_to_bs_82),
			.mem_to_bs_83    (mem_to_bs_83),
			.mem_to_bs_84    (mem_to_bs_84),
			.mem_to_cnu_0    (mem_to_cnu_0),
			.mem_to_cnu_1    (mem_to_cnu_1),
			.mem_to_cnu_2    (mem_to_cnu_2),
			.mem_to_cnu_3    (mem_to_cnu_3),
			.mem_to_cnu_4    (mem_to_cnu_4),
			.mem_to_cnu_5    (mem_to_cnu_5),
			.mem_to_cnu_6    (mem_to_cnu_6),
			.mem_to_cnu_7    (mem_to_cnu_7),
			.mem_to_cnu_8    (mem_to_cnu_8),
			.mem_to_cnu_9    (mem_to_cnu_9),
			.mem_to_cnu_10   (mem_to_cnu_10),
			.mem_to_cnu_11   (mem_to_cnu_11),
			.mem_to_cnu_12   (mem_to_cnu_12),
			.mem_to_cnu_13   (mem_to_cnu_13),
			.mem_to_cnu_14   (mem_to_cnu_14),
			.mem_to_cnu_15   (mem_to_cnu_15),
			.mem_to_cnu_16   (mem_to_cnu_16),
			.mem_to_cnu_17   (mem_to_cnu_17),
			.mem_to_cnu_18   (mem_to_cnu_18),
			.mem_to_cnu_19   (mem_to_cnu_19),
			.mem_to_cnu_20   (mem_to_cnu_20),
			.mem_to_cnu_21   (mem_to_cnu_21),
			.mem_to_cnu_22   (mem_to_cnu_22),
			.mem_to_cnu_23   (mem_to_cnu_23),
			.mem_to_cnu_24   (mem_to_cnu_24),
			.mem_to_cnu_25   (mem_to_cnu_25),
			.mem_to_cnu_26   (mem_to_cnu_26),
			.mem_to_cnu_27   (mem_to_cnu_27),
			.mem_to_cnu_28   (mem_to_cnu_28),
			.mem_to_cnu_29   (mem_to_cnu_29),
			.mem_to_cnu_30   (mem_to_cnu_30),
			.mem_to_cnu_31   (mem_to_cnu_31),
			.mem_to_cnu_32   (mem_to_cnu_32),
			.mem_to_cnu_33   (mem_to_cnu_33),
			.mem_to_cnu_34   (mem_to_cnu_34),
			.mem_to_cnu_35   (mem_to_cnu_35),
			.mem_to_cnu_36   (mem_to_cnu_36),
			.mem_to_cnu_37   (mem_to_cnu_37),
			.mem_to_cnu_38   (mem_to_cnu_38),
			.mem_to_cnu_39   (mem_to_cnu_39),
			.mem_to_cnu_40   (mem_to_cnu_40),
			.mem_to_cnu_41   (mem_to_cnu_41),
			.mem_to_cnu_42   (mem_to_cnu_42),
			.mem_to_cnu_43   (mem_to_cnu_43),
			.mem_to_cnu_44   (mem_to_cnu_44),
			.mem_to_cnu_45   (mem_to_cnu_45),
			.mem_to_cnu_46   (mem_to_cnu_46),
			.mem_to_cnu_47   (mem_to_cnu_47),
			.mem_to_cnu_48   (mem_to_cnu_48),
			.mem_to_cnu_49   (mem_to_cnu_49),
			.mem_to_cnu_50   (mem_to_cnu_50),
			.mem_to_cnu_51   (mem_to_cnu_51),
			.mem_to_cnu_52   (mem_to_cnu_52),
			.mem_to_cnu_53   (mem_to_cnu_53),
			.mem_to_cnu_54   (mem_to_cnu_54),
			.mem_to_cnu_55   (mem_to_cnu_55),
			.mem_to_cnu_56   (mem_to_cnu_56),
			.mem_to_cnu_57   (mem_to_cnu_57),
			.mem_to_cnu_58   (mem_to_cnu_58),
			.mem_to_cnu_59   (mem_to_cnu_59),
			.mem_to_cnu_60   (mem_to_cnu_60),
			.mem_to_cnu_61   (mem_to_cnu_61),
			.mem_to_cnu_62   (mem_to_cnu_62),
			.mem_to_cnu_63   (mem_to_cnu_63),
			.mem_to_cnu_64   (mem_to_cnu_64),
			.mem_to_cnu_65   (mem_to_cnu_65),
			.mem_to_cnu_66   (mem_to_cnu_66),
			.mem_to_cnu_67   (mem_to_cnu_67),
			.mem_to_cnu_68   (mem_to_cnu_68),
			.mem_to_cnu_69   (mem_to_cnu_69),
			.mem_to_cnu_70   (mem_to_cnu_70),
			.mem_to_cnu_71   (mem_to_cnu_71),
			.mem_to_cnu_72   (mem_to_cnu_72),
			.mem_to_cnu_73   (mem_to_cnu_73),
			.mem_to_cnu_74   (mem_to_cnu_74),
			.mem_to_cnu_75   (mem_to_cnu_75),
			.mem_to_cnu_76   (mem_to_cnu_76),
			.mem_to_cnu_77   (mem_to_cnu_77),
			.mem_to_cnu_78   (mem_to_cnu_78),
			.mem_to_cnu_79   (mem_to_cnu_79),
			.mem_to_cnu_80   (mem_to_cnu_80),
			.mem_to_cnu_81   (mem_to_cnu_81),
			.mem_to_cnu_82   (mem_to_cnu_82),
			.mem_to_cnu_83   (mem_to_cnu_83),
			.mem_to_cnu_84   (mem_to_cnu_84),
			.vnu_to_mem_1    (vnu_to_mem_1),
			.vnu_to_mem_1    (vnu_to_mem_1),
			.vnu_to_mem_2    (vnu_to_mem_2),
			.vnu_to_mem_3    (vnu_to_mem_3),
			.vnu_to_mem_4    (vnu_to_mem_4),
			.vnu_to_mem_5    (vnu_to_mem_5),
			.vnu_to_mem_6    (vnu_to_mem_6),
			.vnu_to_mem_7    (vnu_to_mem_7),
			.vnu_to_mem_8    (vnu_to_mem_8),
			.vnu_to_mem_9    (vnu_to_mem_9),
			.vnu_to_mem_10   (vnu_to_mem_10),
			.vnu_to_mem_11   (vnu_to_mem_11),
			.vnu_to_mem_12   (vnu_to_mem_12),
			.vnu_to_mem_13   (vnu_to_mem_13),
			.vnu_to_mem_14   (vnu_to_mem_14),
			.vnu_to_mem_15   (vnu_to_mem_15),
			.vnu_to_mem_16   (vnu_to_mem_16),
			.vnu_to_mem_17   (vnu_to_mem_17),
			.vnu_to_mem_18   (vnu_to_mem_18),
			.vnu_to_mem_19   (vnu_to_mem_19),
			.vnu_to_mem_20   (vnu_to_mem_20),
			.vnu_to_mem_21   (vnu_to_mem_21),
			.vnu_to_mem_22   (vnu_to_mem_22),
			.vnu_to_mem_23   (vnu_to_mem_23),
			.vnu_to_mem_24   (vnu_to_mem_24),
			.vnu_to_mem_25   (vnu_to_mem_25),
			.vnu_to_mem_26   (vnu_to_mem_26),
			.vnu_to_mem_27   (vnu_to_mem_27),
			.vnu_to_mem_28   (vnu_to_mem_28),
			.vnu_to_mem_29   (vnu_to_mem_29),
			.vnu_to_mem_30   (vnu_to_mem_30),
			.vnu_to_mem_31   (vnu_to_mem_31),
			.vnu_to_mem_32   (vnu_to_mem_32),
			.vnu_to_mem_33   (vnu_to_mem_33),
			.vnu_to_mem_34   (vnu_to_mem_34),
			.vnu_to_mem_35   (vnu_to_mem_35),
			.vnu_to_mem_36   (vnu_to_mem_36),
			.vnu_to_mem_37   (vnu_to_mem_37),
			.vnu_to_mem_38   (vnu_to_mem_38),
			.vnu_to_mem_39   (vnu_to_mem_39),
			.vnu_to_mem_40   (vnu_to_mem_40),
			.vnu_to_mem_41   (vnu_to_mem_41),
			.vnu_to_mem_42   (vnu_to_mem_42),
			.vnu_to_mem_43   (vnu_to_mem_43),
			.vnu_to_mem_44   (vnu_to_mem_44),
			.vnu_to_mem_45   (vnu_to_mem_45),
			.vnu_to_mem_46   (vnu_to_mem_46),
			.vnu_to_mem_47   (vnu_to_mem_47),
			.vnu_to_mem_48   (vnu_to_mem_48),
			.vnu_to_mem_49   (vnu_to_mem_49),
			.vnu_to_mem_50   (vnu_to_mem_50),
			.vnu_to_mem_51   (vnu_to_mem_51),
			.vnu_to_mem_52   (vnu_to_mem_52),
			.vnu_to_mem_53   (vnu_to_mem_53),
			.vnu_to_mem_54   (vnu_to_mem_54),
			.vnu_to_mem_55   (vnu_to_mem_55),
			.vnu_to_mem_56   (vnu_to_mem_56),
			.vnu_to_mem_57   (vnu_to_mem_57),
			.vnu_to_mem_58   (vnu_to_mem_58),
			.vnu_to_mem_59   (vnu_to_mem_59),
			.vnu_to_mem_60   (vnu_to_mem_60),
			.vnu_to_mem_61   (vnu_to_mem_61),
			.vnu_to_mem_62   (vnu_to_mem_62),
			.vnu_to_mem_63   (vnu_to_mem_63),
			.vnu_to_mem_64   (vnu_to_mem_64),
			.vnu_to_mem_65   (vnu_to_mem_65),
			.vnu_to_mem_66   (vnu_to_mem_66),
			.vnu_to_mem_67   (vnu_to_mem_67),
			.vnu_to_mem_68   (vnu_to_mem_68),
			.vnu_to_mem_69   (vnu_to_mem_69),
			.vnu_to_mem_70   (vnu_to_mem_70),
			.vnu_to_mem_71   (vnu_to_mem_71),
			.vnu_to_mem_72   (vnu_to_mem_72),
			.vnu_to_mem_73   (vnu_to_mem_73),
			.vnu_to_mem_74   (vnu_to_mem_74),
			.vnu_to_mem_75   (vnu_to_mem_75),
			.vnu_to_mem_76   (vnu_to_mem_76),
			.vnu_to_mem_77   (vnu_to_mem_77),
			.vnu_to_mem_78   (vnu_to_mem_78),
			.vnu_to_mem_79   (vnu_to_mem_79),
			.vnu_to_mem_80   (vnu_to_mem_80),
			.vnu_to_mem_81   (vnu_to_mem_81),
			.vnu_to_mem_82   (vnu_to_mem_82),
			.vnu_to_mem_83   (vnu_to_mem_83),
			.vnu_to_mem_84   (vnu_to_mem_84),
			.cnu_to_mem_0    (cnu_to_mem_0),
			.cnu_to_mem_1    (cnu_to_mem_1),
			.cnu_to_mem_2    (cnu_to_mem_2),
			.cnu_to_mem_3    (cnu_to_mem_3),
			.cnu_to_mem_4    (cnu_to_mem_4),
			.cnu_to_mem_5    (cnu_to_mem_5),
			.cnu_to_mem_6    (cnu_to_mem_6),
			.cnu_to_mem_7    (cnu_to_mem_7),
			.cnu_to_mem_8    (cnu_to_mem_8),
			.cnu_to_mem_9    (cnu_to_mem_9),
			.cnu_to_mem_10   (cnu_to_mem_10),
			.cnu_to_mem_11   (cnu_to_mem_11),
			.cnu_to_mem_12   (cnu_to_mem_12),
			.cnu_to_mem_13   (cnu_to_mem_13),
			.cnu_to_mem_14   (cnu_to_mem_14),
			.cnu_to_mem_15   (cnu_to_mem_15),
			.cnu_to_mem_16   (cnu_to_mem_16),
			.cnu_to_mem_17   (cnu_to_mem_17),
			.cnu_to_mem_18   (cnu_to_mem_18),
			.cnu_to_mem_19   (cnu_to_mem_19),
			.cnu_to_mem_20   (cnu_to_mem_20),
			.cnu_to_mem_21   (cnu_to_mem_21),
			.cnu_to_mem_22   (cnu_to_mem_22),
			.cnu_to_mem_23   (cnu_to_mem_23),
			.cnu_to_mem_24   (cnu_to_mem_24),
			.cnu_to_mem_25   (cnu_to_mem_25),
			.cnu_to_mem_26   (cnu_to_mem_26),
			.cnu_to_mem_27   (cnu_to_mem_27),
			.cnu_to_mem_28   (cnu_to_mem_28),
			.cnu_to_mem_29   (cnu_to_mem_29),
			.cnu_to_mem_30   (cnu_to_mem_30),
			.cnu_to_mem_31   (cnu_to_mem_31),
			.cnu_to_mem_32   (cnu_to_mem_32),
			.cnu_to_mem_33   (cnu_to_mem_33),
			.cnu_to_mem_34   (cnu_to_mem_34),
			.cnu_to_mem_35   (cnu_to_mem_35),
			.cnu_to_mem_36   (cnu_to_mem_36),
			.cnu_to_mem_37   (cnu_to_mem_37),
			.cnu_to_mem_38   (cnu_to_mem_38),
			.cnu_to_mem_39   (cnu_to_mem_39),
			.cnu_to_mem_40   (cnu_to_mem_40),
			.cnu_to_mem_41   (cnu_to_mem_41),
			.cnu_to_mem_42   (cnu_to_mem_42),
			.cnu_to_mem_43   (cnu_to_mem_43),
			.cnu_to_mem_44   (cnu_to_mem_44),
			.cnu_to_mem_45   (cnu_to_mem_45),
			.cnu_to_mem_46   (cnu_to_mem_46),
			.cnu_to_mem_47   (cnu_to_mem_47),
			.cnu_to_mem_48   (cnu_to_mem_48),
			.cnu_to_mem_49   (cnu_to_mem_49),
			.cnu_to_mem_50   (cnu_to_mem_50),
			.cnu_to_mem_51   (cnu_to_mem_51),
			.cnu_to_mem_52   (cnu_to_mem_52),
			.cnu_to_mem_53   (cnu_to_mem_53),
			.cnu_to_mem_54   (cnu_to_mem_54),
			.cnu_to_mem_55   (cnu_to_mem_55),
			.cnu_to_mem_56   (cnu_to_mem_56),
			.cnu_to_mem_57   (cnu_to_mem_57),
			.cnu_to_mem_58   (cnu_to_mem_58),
			.cnu_to_mem_59   (cnu_to_mem_59),
			.cnu_to_mem_60   (cnu_to_mem_60),
			.cnu_to_mem_61   (cnu_to_mem_61),
			.cnu_to_mem_62   (cnu_to_mem_62),
			.cnu_to_mem_63   (cnu_to_mem_63),
			.cnu_to_mem_64   (cnu_to_mem_64),
			.cnu_to_mem_65   (cnu_to_mem_65),
			.cnu_to_mem_66   (cnu_to_mem_66),
			.cnu_to_mem_67   (cnu_to_mem_67),
			.cnu_to_mem_68   (cnu_to_mem_68),
			.cnu_to_mem_69   (cnu_to_mem_69),
			.cnu_to_mem_70   (cnu_to_mem_70),
			.cnu_to_mem_71   (cnu_to_mem_71),
			.cnu_to_mem_72   (cnu_to_mem_72),
			.cnu_to_mem_73   (cnu_to_mem_73),
			.cnu_to_mem_74   (cnu_to_mem_74),
			.cnu_to_mem_75   (cnu_to_mem_75),
			.cnu_to_mem_76   (cnu_to_mem_76),
			.cnu_to_mem_77   (cnu_to_mem_77),
			.cnu_to_mem_78   (cnu_to_mem_78),
			.cnu_to_mem_79   (cnu_to_mem_79),
			.cnu_to_mem_80   (cnu_to_mem_80),
			.cnu_to_mem_81   (cnu_to_mem_81),
			.cnu_to_mem_82   (cnu_to_mem_82),
			.cnu_to_mem_83   (cnu_to_mem_83),
			.cnu_to_mem_84   (cnu_to_mem_84),
			.sched_cmd       (sched_cmd),
			.delay_cmd       (delay_cmd),
			.sync_addr       (sync_addr),
			.layer_status    (layer_status),
			.first_row_chunk (first_row_chunk),
			.we              (we),
			.sys_clk         (sys_clk),
			.rstn            (rstn)
		);

	task init();
		vnu_to_mem_1    <= '0;
		vnu_to_mem_1    <= '0;
		vnu_to_mem_2    <= '0;
		vnu_to_mem_3    <= '0;
		vnu_to_mem_4    <= '0;
		vnu_to_mem_5    <= '0;
		vnu_to_mem_6    <= '0;
		vnu_to_mem_7    <= '0;
		vnu_to_mem_8    <= '0;
		vnu_to_mem_9    <= '0;
		vnu_to_mem_10   <= '0;
		vnu_to_mem_11   <= '0;
		vnu_to_mem_12   <= '0;
		vnu_to_mem_13   <= '0;
		vnu_to_mem_14   <= '0;
		vnu_to_mem_15   <= '0;
		vnu_to_mem_16   <= '0;
		vnu_to_mem_17   <= '0;
		vnu_to_mem_18   <= '0;
		vnu_to_mem_19   <= '0;
		vnu_to_mem_20   <= '0;
		vnu_to_mem_21   <= '0;
		vnu_to_mem_22   <= '0;
		vnu_to_mem_23   <= '0;
		vnu_to_mem_24   <= '0;
		vnu_to_mem_25   <= '0;
		vnu_to_mem_26   <= '0;
		vnu_to_mem_27   <= '0;
		vnu_to_mem_28   <= '0;
		vnu_to_mem_29   <= '0;
		vnu_to_mem_30   <= '0;
		vnu_to_mem_31   <= '0;
		vnu_to_mem_32   <= '0;
		vnu_to_mem_33   <= '0;
		vnu_to_mem_34   <= '0;
		vnu_to_mem_35   <= '0;
		vnu_to_mem_36   <= '0;
		vnu_to_mem_37   <= '0;
		vnu_to_mem_38   <= '0;
		vnu_to_mem_39   <= '0;
		vnu_to_mem_40   <= '0;
		vnu_to_mem_41   <= '0;
		vnu_to_mem_42   <= '0;
		vnu_to_mem_43   <= '0;
		vnu_to_mem_44   <= '0;
		vnu_to_mem_45   <= '0;
		vnu_to_mem_46   <= '0;
		vnu_to_mem_47   <= '0;
		vnu_to_mem_48   <= '0;
		vnu_to_mem_49   <= '0;
		vnu_to_mem_50   <= '0;
		vnu_to_mem_51   <= '0;
		vnu_to_mem_52   <= '0;
		vnu_to_mem_53   <= '0;
		vnu_to_mem_54   <= '0;
		vnu_to_mem_55   <= '0;
		vnu_to_mem_56   <= '0;
		vnu_to_mem_57   <= '0;
		vnu_to_mem_58   <= '0;
		vnu_to_mem_59   <= '0;
		vnu_to_mem_60   <= '0;
		vnu_to_mem_61   <= '0;
		vnu_to_mem_62   <= '0;
		vnu_to_mem_63   <= '0;
		vnu_to_mem_64   <= '0;
		vnu_to_mem_65   <= '0;
		vnu_to_mem_66   <= '0;
		vnu_to_mem_67   <= '0;
		vnu_to_mem_68   <= '0;
		vnu_to_mem_69   <= '0;
		vnu_to_mem_70   <= '0;
		vnu_to_mem_71   <= '0;
		vnu_to_mem_72   <= '0;
		vnu_to_mem_73   <= '0;
		vnu_to_mem_74   <= '0;
		vnu_to_mem_75   <= '0;
		vnu_to_mem_76   <= '0;
		vnu_to_mem_77   <= '0;
		vnu_to_mem_78   <= '0;
		vnu_to_mem_79   <= '0;
		vnu_to_mem_80   <= '0;
		vnu_to_mem_81   <= '0;
		vnu_to_mem_82   <= '0;
		vnu_to_mem_83   <= '0;
		vnu_to_mem_84   <= '0;
		cnu_to_mem_0    <= '0;
		cnu_to_mem_1    <= '0;
		cnu_to_mem_2    <= '0;
		cnu_to_mem_3    <= '0;
		cnu_to_mem_4    <= '0;
		cnu_to_mem_5    <= '0;
		cnu_to_mem_6    <= '0;
		cnu_to_mem_7    <= '0;
		cnu_to_mem_8    <= '0;
		cnu_to_mem_9    <= '0;
		cnu_to_mem_10   <= '0;
		cnu_to_mem_11   <= '0;
		cnu_to_mem_12   <= '0;
		cnu_to_mem_13   <= '0;
		cnu_to_mem_14   <= '0;
		cnu_to_mem_15   <= '0;
		cnu_to_mem_16   <= '0;
		cnu_to_mem_17   <= '0;
		cnu_to_mem_18   <= '0;
		cnu_to_mem_19   <= '0;
		cnu_to_mem_20   <= '0;
		cnu_to_mem_21   <= '0;
		cnu_to_mem_22   <= '0;
		cnu_to_mem_23   <= '0;
		cnu_to_mem_24   <= '0;
		cnu_to_mem_25   <= '0;
		cnu_to_mem_26   <= '0;
		cnu_to_mem_27   <= '0;
		cnu_to_mem_28   <= '0;
		cnu_to_mem_29   <= '0;
		cnu_to_mem_30   <= '0;
		cnu_to_mem_31   <= '0;
		cnu_to_mem_32   <= '0;
		cnu_to_mem_33   <= '0;
		cnu_to_mem_34   <= '0;
		cnu_to_mem_35   <= '0;
		cnu_to_mem_36   <= '0;
		cnu_to_mem_37   <= '0;
		cnu_to_mem_38   <= '0;
		cnu_to_mem_39   <= '0;
		cnu_to_mem_40   <= '0;
		cnu_to_mem_41   <= '0;
		cnu_to_mem_42   <= '0;
		cnu_to_mem_43   <= '0;
		cnu_to_mem_44   <= '0;
		cnu_to_mem_45   <= '0;
		cnu_to_mem_46   <= '0;
		cnu_to_mem_47   <= '0;
		cnu_to_mem_48   <= '0;
		cnu_to_mem_49   <= '0;
		cnu_to_mem_50   <= '0;
		cnu_to_mem_51   <= '0;
		cnu_to_mem_52   <= '0;
		cnu_to_mem_53   <= '0;
		cnu_to_mem_54   <= '0;
		cnu_to_mem_55   <= '0;
		cnu_to_mem_56   <= '0;
		cnu_to_mem_57   <= '0;
		cnu_to_mem_58   <= '0;
		cnu_to_mem_59   <= '0;
		cnu_to_mem_60   <= '0;
		cnu_to_mem_61   <= '0;
		cnu_to_mem_62   <= '0;
		cnu_to_mem_63   <= '0;
		cnu_to_mem_64   <= '0;
		cnu_to_mem_65   <= '0;
		cnu_to_mem_66   <= '0;
		cnu_to_mem_67   <= '0;
		cnu_to_mem_68   <= '0;
		cnu_to_mem_69   <= '0;
		cnu_to_mem_70   <= '0;
		cnu_to_mem_71   <= '0;
		cnu_to_mem_72   <= '0;
		cnu_to_mem_73   <= '0;
		cnu_to_mem_74   <= '0;
		cnu_to_mem_75   <= '0;
		cnu_to_mem_76   <= '0;
		cnu_to_mem_77   <= '0;
		cnu_to_mem_78   <= '0;
		cnu_to_mem_79   <= '0;
		cnu_to_mem_80   <= '0;
		cnu_to_mem_81   <= '0;
		cnu_to_mem_82   <= '0;
		cnu_to_mem_83   <= '0;
		cnu_to_mem_84   <= '0;
		sched_cmd       <= '0;
		delay_cmd       <= '0;
		sync_addr       <= '0;
		layer_status    <= '0;
		first_row_chunk <= '0;
		we              <= '0;
		sys_clk         <= '0;
		rstn            <= '0;
	endtask

	task drive(int iter);
		for(int it = 0; it < iter; it++) begin
			vnu_to_mem_1    <= '0;
			vnu_to_mem_1    <= '0;
			vnu_to_mem_2    <= '0;
			vnu_to_mem_3    <= '0;
			vnu_to_mem_4    <= '0;
			vnu_to_mem_5    <= '0;
			vnu_to_mem_6    <= '0;
			vnu_to_mem_7    <= '0;
			vnu_to_mem_8    <= '0;
			vnu_to_mem_9    <= '0;
			vnu_to_mem_10   <= '0;
			vnu_to_mem_11   <= '0;
			vnu_to_mem_12   <= '0;
			vnu_to_mem_13   <= '0;
			vnu_to_mem_14   <= '0;
			vnu_to_mem_15   <= '0;
			vnu_to_mem_16   <= '0;
			vnu_to_mem_17   <= '0;
			vnu_to_mem_18   <= '0;
			vnu_to_mem_19   <= '0;
			vnu_to_mem_20   <= '0;
			vnu_to_mem_21   <= '0;
			vnu_to_mem_22   <= '0;
			vnu_to_mem_23   <= '0;
			vnu_to_mem_24   <= '0;
			vnu_to_mem_25   <= '0;
			vnu_to_mem_26   <= '0;
			vnu_to_mem_27   <= '0;
			vnu_to_mem_28   <= '0;
			vnu_to_mem_29   <= '0;
			vnu_to_mem_30   <= '0;
			vnu_to_mem_31   <= '0;
			vnu_to_mem_32   <= '0;
			vnu_to_mem_33   <= '0;
			vnu_to_mem_34   <= '0;
			vnu_to_mem_35   <= '0;
			vnu_to_mem_36   <= '0;
			vnu_to_mem_37   <= '0;
			vnu_to_mem_38   <= '0;
			vnu_to_mem_39   <= '0;
			vnu_to_mem_40   <= '0;
			vnu_to_mem_41   <= '0;
			vnu_to_mem_42   <= '0;
			vnu_to_mem_43   <= '0;
			vnu_to_mem_44   <= '0;
			vnu_to_mem_45   <= '0;
			vnu_to_mem_46   <= '0;
			vnu_to_mem_47   <= '0;
			vnu_to_mem_48   <= '0;
			vnu_to_mem_49   <= '0;
			vnu_to_mem_50   <= '0;
			vnu_to_mem_51   <= '0;
			vnu_to_mem_52   <= '0;
			vnu_to_mem_53   <= '0;
			vnu_to_mem_54   <= '0;
			vnu_to_mem_55   <= '0;
			vnu_to_mem_56   <= '0;
			vnu_to_mem_57   <= '0;
			vnu_to_mem_58   <= '0;
			vnu_to_mem_59   <= '0;
			vnu_to_mem_60   <= '0;
			vnu_to_mem_61   <= '0;
			vnu_to_mem_62   <= '0;
			vnu_to_mem_63   <= '0;
			vnu_to_mem_64   <= '0;
			vnu_to_mem_65   <= '0;
			vnu_to_mem_66   <= '0;
			vnu_to_mem_67   <= '0;
			vnu_to_mem_68   <= '0;
			vnu_to_mem_69   <= '0;
			vnu_to_mem_70   <= '0;
			vnu_to_mem_71   <= '0;
			vnu_to_mem_72   <= '0;
			vnu_to_mem_73   <= '0;
			vnu_to_mem_74   <= '0;
			vnu_to_mem_75   <= '0;
			vnu_to_mem_76   <= '0;
			vnu_to_mem_77   <= '0;
			vnu_to_mem_78   <= '0;
			vnu_to_mem_79   <= '0;
			vnu_to_mem_80   <= '0;
			vnu_to_mem_81   <= '0;
			vnu_to_mem_82   <= '0;
			vnu_to_mem_83   <= '0;
			vnu_to_mem_84   <= '0;
			cnu_to_mem_0    <= '0;
			cnu_to_mem_1    <= '0;
			cnu_to_mem_2    <= '0;
			cnu_to_mem_3    <= '0;
			cnu_to_mem_4    <= '0;
			cnu_to_mem_5    <= '0;
			cnu_to_mem_6    <= '0;
			cnu_to_mem_7    <= '0;
			cnu_to_mem_8    <= '0;
			cnu_to_mem_9    <= '0;
			cnu_to_mem_10   <= '0;
			cnu_to_mem_11   <= '0;
			cnu_to_mem_12   <= '0;
			cnu_to_mem_13   <= '0;
			cnu_to_mem_14   <= '0;
			cnu_to_mem_15   <= '0;
			cnu_to_mem_16   <= '0;
			cnu_to_mem_17   <= '0;
			cnu_to_mem_18   <= '0;
			cnu_to_mem_19   <= '0;
			cnu_to_mem_20   <= '0;
			cnu_to_mem_21   <= '0;
			cnu_to_mem_22   <= '0;
			cnu_to_mem_23   <= '0;
			cnu_to_mem_24   <= '0;
			cnu_to_mem_25   <= '0;
			cnu_to_mem_26   <= '0;
			cnu_to_mem_27   <= '0;
			cnu_to_mem_28   <= '0;
			cnu_to_mem_29   <= '0;
			cnu_to_mem_30   <= '0;
			cnu_to_mem_31   <= '0;
			cnu_to_mem_32   <= '0;
			cnu_to_mem_33   <= '0;
			cnu_to_mem_34   <= '0;
			cnu_to_mem_35   <= '0;
			cnu_to_mem_36   <= '0;
			cnu_to_mem_37   <= '0;
			cnu_to_mem_38   <= '0;
			cnu_to_mem_39   <= '0;
			cnu_to_mem_40   <= '0;
			cnu_to_mem_41   <= '0;
			cnu_to_mem_42   <= '0;
			cnu_to_mem_43   <= '0;
			cnu_to_mem_44   <= '0;
			cnu_to_mem_45   <= '0;
			cnu_to_mem_46   <= '0;
			cnu_to_mem_47   <= '0;
			cnu_to_mem_48   <= '0;
			cnu_to_mem_49   <= '0;
			cnu_to_mem_50   <= '0;
			cnu_to_mem_51   <= '0;
			cnu_to_mem_52   <= '0;
			cnu_to_mem_53   <= '0;
			cnu_to_mem_54   <= '0;
			cnu_to_mem_55   <= '0;
			cnu_to_mem_56   <= '0;
			cnu_to_mem_57   <= '0;
			cnu_to_mem_58   <= '0;
			cnu_to_mem_59   <= '0;
			cnu_to_mem_60   <= '0;
			cnu_to_mem_61   <= '0;
			cnu_to_mem_62   <= '0;
			cnu_to_mem_63   <= '0;
			cnu_to_mem_64   <= '0;
			cnu_to_mem_65   <= '0;
			cnu_to_mem_66   <= '0;
			cnu_to_mem_67   <= '0;
			cnu_to_mem_68   <= '0;
			cnu_to_mem_69   <= '0;
			cnu_to_mem_70   <= '0;
			cnu_to_mem_71   <= '0;
			cnu_to_mem_72   <= '0;
			cnu_to_mem_73   <= '0;
			cnu_to_mem_74   <= '0;
			cnu_to_mem_75   <= '0;
			cnu_to_mem_76   <= '0;
			cnu_to_mem_77   <= '0;
			cnu_to_mem_78   <= '0;
			cnu_to_mem_79   <= '0;
			cnu_to_mem_80   <= '0;
			cnu_to_mem_81   <= '0;
			cnu_to_mem_82   <= '0;
			cnu_to_mem_83   <= '0;
			cnu_to_mem_84   <= '0;
			sched_cmd       <= '0;
			delay_cmd       <= '0;
			sync_addr       <= '0;
			layer_status    <= '0;
			first_row_chunk <= '0;
			we              <= '0;
			sys_clk         <= '0;
			rstn            <= '0;
			@(posedge clk);
		end
	endtask

	initial begin
		// do something

		init();
		repeat(10)@(posedge clk);

		drive(20);

		repeat(10)@(posedge clk);
		$finish;
	end

	// dump wave
	initial begin
		$display("random seed : %0d", $unsigned($get_initial_random_seed()));
		if ( $test$plusargs("fsdb") ) begin
			$fsdbDumpfile("tb_mem_subsystem_top.fsdb");
			$fsdbDumpvars(0, "tb_mem_subsystem_top", "+mda", "+functions");
		end
	end

endmodule