`include "define.vh"

`ifdef SCHED_4_6
module ram_pageAlign_interface_submatrix_2#(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 85,
	parameter LAYER_NUM = 3
) (
	output wire [QUAN_SIZE-1:0] msg_out_0,
	output wire [QUAN_SIZE-1:0] msg_out_1,
	output wire [QUAN_SIZE-1:0] msg_out_2,
	output wire [QUAN_SIZE-1:0] msg_out_3,
	output wire [QUAN_SIZE-1:0] msg_out_4,
	output wire [QUAN_SIZE-1:0] msg_out_5,
	output wire [QUAN_SIZE-1:0] msg_out_6,
	output wire [QUAN_SIZE-1:0] msg_out_7,
	output wire [QUAN_SIZE-1:0] msg_out_8,
	output wire [QUAN_SIZE-1:0] msg_out_9,
	output wire [QUAN_SIZE-1:0] msg_out_10,
	output wire [QUAN_SIZE-1:0] msg_out_11,
	output wire [QUAN_SIZE-1:0] msg_out_12,
	output wire [QUAN_SIZE-1:0] msg_out_13,
	output wire [QUAN_SIZE-1:0] msg_out_14,
	output wire [QUAN_SIZE-1:0] msg_out_15,
	output wire [QUAN_SIZE-1:0] msg_out_16,
	output wire [QUAN_SIZE-1:0] msg_out_17,
	output wire [QUAN_SIZE-1:0] msg_out_18,
	output wire [QUAN_SIZE-1:0] msg_out_19,
	output wire [QUAN_SIZE-1:0] msg_out_20,
	output wire [QUAN_SIZE-1:0] msg_out_21,
	output wire [QUAN_SIZE-1:0] msg_out_22,
	output wire [QUAN_SIZE-1:0] msg_out_23,
	output wire [QUAN_SIZE-1:0] msg_out_24,
	output wire [QUAN_SIZE-1:0] msg_out_25,
	output wire [QUAN_SIZE-1:0] msg_out_26,
	output wire [QUAN_SIZE-1:0] msg_out_27,
	output wire [QUAN_SIZE-1:0] msg_out_28,
	output wire [QUAN_SIZE-1:0] msg_out_29,
	output wire [QUAN_SIZE-1:0] msg_out_30,
	output wire [QUAN_SIZE-1:0] msg_out_31,
	output wire [QUAN_SIZE-1:0] msg_out_32,
	output wire [QUAN_SIZE-1:0] msg_out_33,
	output wire [QUAN_SIZE-1:0] msg_out_34,
	output wire [QUAN_SIZE-1:0] msg_out_35,
	output wire [QUAN_SIZE-1:0] msg_out_36,
	output wire [QUAN_SIZE-1:0] msg_out_37,
	output wire [QUAN_SIZE-1:0] msg_out_38,
	output wire [QUAN_SIZE-1:0] msg_out_39,
	output wire [QUAN_SIZE-1:0] msg_out_40,
	output wire [QUAN_SIZE-1:0] msg_out_41,
	output wire [QUAN_SIZE-1:0] msg_out_42,
	output wire [QUAN_SIZE-1:0] msg_out_43,
	output wire [QUAN_SIZE-1:0] msg_out_44,
	output wire [QUAN_SIZE-1:0] msg_out_45,
	output wire [QUAN_SIZE-1:0] msg_out_46,
	output wire [QUAN_SIZE-1:0] msg_out_47,
	output wire [QUAN_SIZE-1:0] msg_out_48,
	output wire [QUAN_SIZE-1:0] msg_out_49,
	output wire [QUAN_SIZE-1:0] msg_out_50,
	output wire [QUAN_SIZE-1:0] msg_out_51,
	output wire [QUAN_SIZE-1:0] msg_out_52,
	output wire [QUAN_SIZE-1:0] msg_out_53,
	output wire [QUAN_SIZE-1:0] msg_out_54,
	output wire [QUAN_SIZE-1:0] msg_out_55,
	output wire [QUAN_SIZE-1:0] msg_out_56,
	output wire [QUAN_SIZE-1:0] msg_out_57,
	output wire [QUAN_SIZE-1:0] msg_out_58,
	output wire [QUAN_SIZE-1:0] msg_out_59,
	output wire [QUAN_SIZE-1:0] msg_out_60,
	output wire [QUAN_SIZE-1:0] msg_out_61,
	output wire [QUAN_SIZE-1:0] msg_out_62,
	output wire [QUAN_SIZE-1:0] msg_out_63,
	output wire [QUAN_SIZE-1:0] msg_out_64,
	output wire [QUAN_SIZE-1:0] msg_out_65,
	output wire [QUAN_SIZE-1:0] msg_out_66,
	output wire [QUAN_SIZE-1:0] msg_out_67,
	output wire [QUAN_SIZE-1:0] msg_out_68,
	output wire [QUAN_SIZE-1:0] msg_out_69,
	output wire [QUAN_SIZE-1:0] msg_out_70,
	output wire [QUAN_SIZE-1:0] msg_out_71,
	output wire [QUAN_SIZE-1:0] msg_out_72,
	output wire [QUAN_SIZE-1:0] msg_out_73,
	output wire [QUAN_SIZE-1:0] msg_out_74,
	output wire [QUAN_SIZE-1:0] msg_out_75,
	output wire [QUAN_SIZE-1:0] msg_out_76,
	output wire [QUAN_SIZE-1:0] msg_out_77,
	output wire [QUAN_SIZE-1:0] msg_out_78,
	output wire [QUAN_SIZE-1:0] msg_out_79,
	output wire [QUAN_SIZE-1:0] msg_out_80,
	output wire [QUAN_SIZE-1:0] msg_out_81,
	output wire [QUAN_SIZE-1:0] msg_out_82,
	output wire [QUAN_SIZE-1:0] msg_out_83,
	output wire [QUAN_SIZE-1:0] msg_out_84,

	input wire [QUAN_SIZE-1:0] msg_in_0,
	input wire [QUAN_SIZE-1:0] msg_in_1,
	input wire [QUAN_SIZE-1:0] msg_in_2,
	input wire [QUAN_SIZE-1:0] msg_in_3,
	input wire [QUAN_SIZE-1:0] msg_in_4,
	input wire [QUAN_SIZE-1:0] msg_in_5,
	input wire [QUAN_SIZE-1:0] msg_in_6,
	input wire [QUAN_SIZE-1:0] msg_in_7,
	input wire [QUAN_SIZE-1:0] msg_in_8,
	input wire [QUAN_SIZE-1:0] msg_in_9,
	input wire [QUAN_SIZE-1:0] msg_in_10,
	input wire [QUAN_SIZE-1:0] msg_in_11,
	input wire [QUAN_SIZE-1:0] msg_in_12,
	input wire [QUAN_SIZE-1:0] msg_in_13,
	input wire [QUAN_SIZE-1:0] msg_in_14,
	input wire [QUAN_SIZE-1:0] msg_in_15,
	input wire [QUAN_SIZE-1:0] msg_in_16,
	input wire [QUAN_SIZE-1:0] msg_in_17,
	input wire [QUAN_SIZE-1:0] msg_in_18,
	input wire [QUAN_SIZE-1:0] msg_in_19,
	input wire [QUAN_SIZE-1:0] msg_in_20,
	input wire [QUAN_SIZE-1:0] msg_in_21,
	input wire [QUAN_SIZE-1:0] msg_in_22,
	input wire [QUAN_SIZE-1:0] msg_in_23,
	input wire [QUAN_SIZE-1:0] msg_in_24,
	input wire [QUAN_SIZE-1:0] msg_in_25,
	input wire [QUAN_SIZE-1:0] msg_in_26,
	input wire [QUAN_SIZE-1:0] msg_in_27,
	input wire [QUAN_SIZE-1:0] msg_in_28,
	input wire [QUAN_SIZE-1:0] msg_in_29,
	input wire [QUAN_SIZE-1:0] msg_in_30,
	input wire [QUAN_SIZE-1:0] msg_in_31,
	input wire [QUAN_SIZE-1:0] msg_in_32,
	input wire [QUAN_SIZE-1:0] msg_in_33,
	input wire [QUAN_SIZE-1:0] msg_in_34,
	input wire [QUAN_SIZE-1:0] msg_in_35,
	input wire [QUAN_SIZE-1:0] msg_in_36,
	input wire [QUAN_SIZE-1:0] msg_in_37,
	input wire [QUAN_SIZE-1:0] msg_in_38,
	input wire [QUAN_SIZE-1:0] msg_in_39,
	input wire [QUAN_SIZE-1:0] msg_in_40,
	input wire [QUAN_SIZE-1:0] msg_in_41,
	input wire [QUAN_SIZE-1:0] msg_in_42,
	input wire [QUAN_SIZE-1:0] msg_in_43,
	input wire [QUAN_SIZE-1:0] msg_in_44,
	input wire [QUAN_SIZE-1:0] msg_in_45,
	input wire [QUAN_SIZE-1:0] msg_in_46,
	input wire [QUAN_SIZE-1:0] msg_in_47,
	input wire [QUAN_SIZE-1:0] msg_in_48,
	input wire [QUAN_SIZE-1:0] msg_in_49,
	input wire [QUAN_SIZE-1:0] msg_in_50,
	input wire [QUAN_SIZE-1:0] msg_in_51,
	input wire [QUAN_SIZE-1:0] msg_in_52,
	input wire [QUAN_SIZE-1:0] msg_in_53,
	input wire [QUAN_SIZE-1:0] msg_in_54,
	input wire [QUAN_SIZE-1:0] msg_in_55,
	input wire [QUAN_SIZE-1:0] msg_in_56,
	input wire [QUAN_SIZE-1:0] msg_in_57,
	input wire [QUAN_SIZE-1:0] msg_in_58,
	input wire [QUAN_SIZE-1:0] msg_in_59,
	input wire [QUAN_SIZE-1:0] msg_in_60,
	input wire [QUAN_SIZE-1:0] msg_in_61,
	input wire [QUAN_SIZE-1:0] msg_in_62,
	input wire [QUAN_SIZE-1:0] msg_in_63,
	input wire [QUAN_SIZE-1:0] msg_in_64,
	input wire [QUAN_SIZE-1:0] msg_in_65,
	input wire [QUAN_SIZE-1:0] msg_in_66,
	input wire [QUAN_SIZE-1:0] msg_in_67,
	input wire [QUAN_SIZE-1:0] msg_in_68,
	input wire [QUAN_SIZE-1:0] msg_in_69,
	input wire [QUAN_SIZE-1:0] msg_in_70,
	input wire [QUAN_SIZE-1:0] msg_in_71,
	input wire [QUAN_SIZE-1:0] msg_in_72,
	input wire [QUAN_SIZE-1:0] msg_in_73,
	input wire [QUAN_SIZE-1:0] msg_in_74,
	input wire [QUAN_SIZE-1:0] msg_in_75,
	input wire [QUAN_SIZE-1:0] msg_in_76,
	input wire [QUAN_SIZE-1:0] msg_in_77,
	input wire [QUAN_SIZE-1:0] msg_in_78,
	input wire [QUAN_SIZE-1:0] msg_in_79,
	input wire [QUAN_SIZE-1:0] msg_in_80,
	input wire [QUAN_SIZE-1:0] msg_in_81,
	input wire [QUAN_SIZE-1:0] msg_in_82,
	input wire [QUAN_SIZE-1:0] msg_in_83,
	input wire [QUAN_SIZE-1:0] msg_in_84,

	input wire [LAYER_NUM-1:0] layer_status,
	input wire first_row_chunk,
	input wire sys_clk,
	input wire rstn
);

/////////////////////////////////////////////////////////////////////////////////////////////
// Main structure of Page Alignment Mechanism
wire [1:0] circular_delay_cmd_3_2;
assign circular_delay_cmd_3_2 = ((layer_status[0] == 1'b1 || layer_status[1] == 1'b1) && first_row_chunk == 1'b1) ? 2'b10 : (layer_status[2] == 1'b1) ? 2'b01 : 2'b00;
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u21 (.align_out (msg_out_21), .align_target_in (msg_in_21), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u22 (.align_out (msg_out_22), .align_target_in (msg_in_22), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u23 (.align_out (msg_out_23), .align_target_in (msg_in_23), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u24 (.align_out (msg_out_24), .align_target_in (msg_in_24), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u25 (.align_out (msg_out_25), .align_target_in (msg_in_25), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u26 (.align_out (msg_out_26), .align_target_in (msg_in_26), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u27 (.align_out (msg_out_27), .align_target_in (msg_in_27), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u28 (.align_out (msg_out_28), .align_target_in (msg_in_28), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u29 (.align_out (msg_out_29), .align_target_in (msg_in_29), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u60 (.align_out (msg_out_60), .align_target_in (msg_in_60), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u61 (.align_out (msg_out_61), .align_target_in (msg_in_61), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u62 (.align_out (msg_out_62), .align_target_in (msg_in_62), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u63 (.align_out (msg_out_63), .align_target_in (msg_in_63), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u64 (.align_out (msg_out_64), .align_target_in (msg_in_64), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u65 (.align_out (msg_out_65), .align_target_in (msg_in_65), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u66 (.align_out (msg_out_66), .align_target_in (msg_in_66), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u67 (.align_out (msg_out_67), .align_target_in (msg_in_67), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u68 (.align_out (msg_out_68), .align_target_in (msg_in_68), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u69 (.align_out (msg_out_69), .align_target_in (msg_in_69), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u70 (.align_out (msg_out_70), .align_target_in (msg_in_70), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u71 (.align_out (msg_out_71), .align_target_in (msg_in_71), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u72 (.align_out (msg_out_72), .align_target_in (msg_in_72), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u73 (.align_out (msg_out_73), .align_target_in (msg_in_73), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u74 (.align_out (msg_out_74), .align_target_in (msg_in_74), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u75 (.align_out (msg_out_75), .align_target_in (msg_in_75), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u76 (.align_out (msg_out_76), .align_target_in (msg_in_76), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u77 (.align_out (msg_out_77), .align_target_in (msg_in_77), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u78 (.align_out (msg_out_78), .align_target_in (msg_in_78), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u79 (.align_out (msg_out_79), .align_target_in (msg_in_79), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u80 (.align_out (msg_out_80), .align_target_in (msg_in_80), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u81 (.align_out (msg_out_81), .align_target_in (msg_in_81), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u82 (.align_out (msg_out_82), .align_target_in (msg_in_82), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u83 (.align_out (msg_out_83), .align_target_in (msg_in_83), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u84 (.align_out (msg_out_84), .align_target_in (msg_in_84), .delay_cmd(circular_delay_cmd_3_2), .sys_clk(sys_clk), .rstn(rstn));
wire [1:0] circular_delay_cmd_5_0;
assign circular_delay_cmd_5_0 = (layer_status[0] == 1'b1 && first_row_chunk == 1'b1) ? 2'b10 : (layer_status[1] == 1'b1 || layer_status[2] == 1'b1) ? 2'b01 : 2'b00;
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u9 (.align_out (msg_out_9), .align_target_in (msg_in_9), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u10 (.align_out (msg_out_10), .align_target_in (msg_in_10), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u11 (.align_out (msg_out_11), .align_target_in (msg_in_11), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u12 (.align_out (msg_out_12), .align_target_in (msg_in_12), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u13 (.align_out (msg_out_13), .align_target_in (msg_in_13), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u14 (.align_out (msg_out_14), .align_target_in (msg_in_14), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u15 (.align_out (msg_out_15), .align_target_in (msg_in_15), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u16 (.align_out (msg_out_16), .align_target_in (msg_in_16), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u17 (.align_out (msg_out_17), .align_target_in (msg_in_17), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u18 (.align_out (msg_out_18), .align_target_in (msg_in_18), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u19 (.align_out (msg_out_19), .align_target_in (msg_in_19), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u20 (.align_out (msg_out_20), .align_target_in (msg_in_20), .delay_cmd(circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u0(.align_out(msg_out_0), .align_target_in (msg_in_0), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u1(.align_out(msg_out_1), .align_target_in (msg_in_1), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u2(.align_out(msg_out_2), .align_target_in (msg_in_2), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u3(.align_out(msg_out_3), .align_target_in (msg_in_3), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u4(.align_out(msg_out_4), .align_target_in (msg_in_4), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u5(.align_out(msg_out_5), .align_target_in (msg_in_5), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u6(.align_out(msg_out_6), .align_target_in (msg_in_6), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u7(.align_out(msg_out_7), .align_target_in (msg_in_7), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u8(.align_out(msg_out_8), .align_target_in (msg_in_8), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u30 (.align_out (msg_out_30), .align_target_in (msg_in_30), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u31 (.align_out (msg_out_31), .align_target_in (msg_in_31), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u32 (.align_out (msg_out_32), .align_target_in (msg_in_32), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u33 (.align_out (msg_out_33), .align_target_in (msg_in_33), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u34 (.align_out (msg_out_34), .align_target_in (msg_in_34), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u35 (.align_out (msg_out_35), .align_target_in (msg_in_35), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u36 (.align_out (msg_out_36), .align_target_in (msg_in_36), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u37 (.align_out (msg_out_37), .align_target_in (msg_in_37), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u38 (.align_out (msg_out_38), .align_target_in (msg_in_38), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u39 (.align_out (msg_out_39), .align_target_in (msg_in_39), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u40 (.align_out (msg_out_40), .align_target_in (msg_in_40), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u41 (.align_out (msg_out_41), .align_target_in (msg_in_41), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u42 (.align_out (msg_out_42), .align_target_in (msg_in_42), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u43 (.align_out (msg_out_43), .align_target_in (msg_in_43), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u44 (.align_out (msg_out_44), .align_target_in (msg_in_44), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u45 (.align_out (msg_out_45), .align_target_in (msg_in_45), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u46 (.align_out (msg_out_46), .align_target_in (msg_in_46), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u47 (.align_out (msg_out_47), .align_target_in (msg_in_47), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u48 (.align_out (msg_out_48), .align_target_in (msg_in_48), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u49 (.align_out (msg_out_49), .align_target_in (msg_in_49), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u50 (.align_out (msg_out_50), .align_target_in (msg_in_50), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u51 (.align_out (msg_out_51), .align_target_in (msg_in_51), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u52 (.align_out (msg_out_52), .align_target_in (msg_in_52), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u53 (.align_out (msg_out_53), .align_target_in (msg_in_53), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u54 (.align_out (msg_out_54), .align_target_in (msg_in_54), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u55 (.align_out (msg_out_55), .align_target_in (msg_in_55), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u56 (.align_out (msg_out_56), .align_target_in (msg_in_56), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u57 (.align_out (msg_out_57), .align_target_in (msg_in_57), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u58 (.align_out (msg_out_58), .align_target_in (msg_in_58), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u59 (.align_out (msg_out_59), .align_target_in (msg_in_59), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
/////////////////////////////////////////////////////////////////////////////////////////////
endmodule
`endif