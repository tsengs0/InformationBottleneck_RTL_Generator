`timescale 1ns / 1ps
`include "define.vh"

module entire_decoder_tb;

// FSM steps for Sys.FSMs
localparam [3:0] INIT_LOAD     = 4'b0000;
localparam [3:0] LLR_FETCH     = 4'b0001;  
localparam [3:0] LLR_FETCH_OUT = 4'b0010;
localparam [3:0] CNU_PIPE      = 4'b0011;
localparam [3:0] CNU_OUT       = 4'b0100;
localparam [3:0] P2P_C         = 4'b0101;
localparam [3:0] P2P_C_OUT     = 4'b0110;
localparam [3:0] VNU_PIPE      = 4'b0111;
localparam [3:0] VNU_OUT       = 4'b1000;
localparam [3:0] P2P_V         = 4'b1001;
localparam [3:0] P2P_V_OUT     = 4'b1010;

//////////////////////////////////////////////////////////////////////////////////////////////////////
// Memory System

// Memory System - Output
/*Check Node*/
wire [CN_RD_BW-1:0] cn_iter0_m0_portA_dout;
wire [CN_RD_BW-1:0] cn_iter0_m0_portB_dout;
wire [CN_RD_BW-1:0] cn_iter0_m1_portA_dout;
wire [CN_RD_BW-1:0] cn_iter0_m1_portB_dout;
wire [CN_RD_BW-1:0] cn_iter0_m2_portA_dout;
wire [CN_RD_BW-1:0] cn_iter0_m2_portB_dout;
wire [CN_RD_BW-1:0] cn_iter0_m3_portA_dout;
wire [CN_RD_BW-1:0] cn_iter0_m3_portB_dout;
wire [CN_RD_BW-1:0] cn_iter1_m0_portA_dout;
wire [CN_RD_BW-1:0] cn_iter1_m0_portB_dout;
wire [CN_RD_BW-1:0] cn_iter1_m1_portA_dout;
wire [CN_RD_BW-1:0] cn_iter1_m1_portB_dout;
wire [CN_RD_BW-1:0] cn_iter1_m2_portA_dout;
wire [CN_RD_BW-1:0] cn_iter1_m2_portB_dout;
wire [CN_RD_BW-1:0] cn_iter1_m3_portA_dout;
wire [CN_RD_BW-1:0] cn_iter1_m3_portB_dout;
/*Variable Node*/
wire [VN_RD_BW-1:0] vn_iter0_m0_portA_dout;
wire [VN_RD_BW-1:0] vn_iter0_m0_portB_dout;
wire [VN_RD_BW-1:0] vn_iter0_m1_portA_dout;
wire [VN_RD_BW-1:0] vn_iter0_m1_portB_dout;
wire [VN_RD_BW-1:0] vn_iter1_m0_portA_dout;
wire [VN_RD_BW-1:0] vn_iter1_m0_portB_dout;
wire [VN_RD_BW-1:0] vn_iter1_m1_portA_dout;
wire [VN_RD_BW-1:0] vn_iter1_m1_portB_dout;
/*Decision Node*/
wire [DN_RD_BW-1:0] dn_iter0_m2_portA_dout;
wire [DN_RD_BW-1:0] dn_iter0_m2_portB_dout;
wire [DN_RD_BW-1:0] dn_iter1_m2_portA_dout;
wire [DN_RD_BW-1:0] dn_iter1_m2_portB_dout;


// Memory System - Ouput of Mux
/*Check Node*/
wire [CN_RD_BW-1:0] cn_portA_dout [0:`IB_CNU_DECOMP_funNum-1];
wire [CN_RD_BW-1:0] cn_portB_dout [0:`IB_CNU_DECOMP_funNum-1];
/*Variable Node*/
wire [VN_RD_BW-1:0] vn_portA_dout [0:`IB_VNU_DECOMP_funNum-1];
wire [VN_RD_BW-1:0] vn_portB_dout [0:`IB_VNU_DECOMP_funNum-1];
/*Decision Node*/
wire [DN_RD_BW-1:0] dn_portA_dout;
wire [DN_RD_BW-1:0] dn_portB_dout;

// Memory Latch - Output
/*Check Node*/
wire [ROM_RD_BW-1:0] cn_latch_outA [0:`IB_CNU_DECOMP_funNum-1];
wire [ROM_RD_BW-1:0] cn_latch_outB [0:`IB_CNU_DECOMP_funNum-1];
wire [ROM_ADDR_BW-1:0] cn_rom_read_addrA [0:`IB_CNU_DECOMP_funNum-1];
wire [ROM_ADDR_BW-1:0] cn_rom_read_addrB [0:`IB_CNU_DECOMP_funNum-1];
/*Variable Node*/
wire [ROM_RD_BW-1:0]   vn_latch_outA [0:`IB_VNU_DECOMP_funNum-1];
wire [ROM_RD_BW-1:0]   vn_latch_outB [0:`IB_VNU_DECOMP_funNum-1];
wire [ROM_ADDR_BW-1:0] vn_rom_read_addrA [0:`IB_VNU_DECOMP_funNum-1];
wire [ROM_ADDR_BW-1:0] vn_rom_read_addrB [0:`IB_VNU_DECOMP_funNum-1];
/*Decision Node*/
wire [ROM_RD_BW-1:0]   dn_latch_outA;
wire [ROM_RD_BW-1:0]   dn_latch_outB;
wire [ROM_ADDR_BW-1:0] dn_rom_read_addrA;
wire [ROM_ADDR_BW-1:0] dn_rom_read_addrB;

// IB-RAM Write Page Address Counter - Output
wire [PAGE_ADDR_BW-1:0] cn_wr_page_addr [0:`IB_CNU_DECOMP_funNum-1];
wire [PAGE_ADDR_BW-1:0] vn_wr_page_addr [0:`IB_VNU_DECOMP_funNum-1];
wire [PAGE_ADDR_BW-1:0] dn_wr_page_addr;
//////////////////////////////////////////////////////////////////////////////////////////////////////
// FSM steps for Write.FSMs
localparam IDLE       = 3'b000;
localparam ROM_FETCH0 = 3'b001; // only for the first write or non-pipeline fashion
localparam RAM_LOAD0  = 3'b010;
localparam RAM_LOAD1  = 3'b011;
localparam FINISH     = 3'b100;

localparam INTER_FRAME_LEVEL = 2;
localparam simulate_iteration = 10; // only simulating until 9th iterations
localparam simulate_codewords = 5; // only simulating until 4th codeword deconding process
localparam iter_cnt_bitwidth = $clog2(simulate_iteration);
localparam codeword_cnt_bitwidth = $clog2(simulate_codewords);
reg [iter_cnt_bitwidth-1:0] iter_cnt;
reg [codeword_cnt_bitwidth-1:0] codeword_cnt;
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Global Simulation Nets
reg cn_write_clk, vn_write_clk, dn_write_clk;
logic [`IB_CNU_DECOMP_funNum-1:0] cn_iter_switch;
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Nets of Sys.FSMs
wire [INTER_FRAME_LEVEL-1:0] llr_fetch;
wire [INTER_FRAME_LEVEL-1:0] v2c_src;
wire [INTER_FRAME_LEVEL-1:0] v2c_msg_en;
wire [`IB_CNU_DECOMP_funNum-1:0] cnu_rd [0:INTER_FRAME_LEVEL-1];
wire [INTER_FRAME_LEVEL-1:0] c2v_msg_en;
wire [`IB_VNU_DECOMP_funNum-1:0] vnu_rd [0:INTER_FRAME_LEVEL-1];
wire dnu_rd [0:INTER_FRAME_LEVEL-1];
wire [INTER_FRAME_LEVEL-1:0] c2v_load;
wire [INTER_FRAME_LEVEL-1:0] v2c_load;
wire [INTER_FRAME_LEVEL-1:0] de_frame_start;
wire [INTER_FRAME_LEVEL-1:0] inter_frame_en;
wire [3:0] sys_fsm_state [0:INTER_FRAME_LEVEL-1];
reg [INTER_FRAME_LEVEL-1:0] fsm_en;
/*Obsoleted*///wire [`IB_CNU_DECOMP_funNum-1:0] fsm_cn_ram_re [0:INTER_FRAME_LEVEL-1];
/*Obsoleted*///wire [`IB_VNU_DECOMP_funNum-1:0] fsm_vn_ram_re [0:INTER_FRAME_LEVEL-1];
/*Obsoleted*///wire [INTER_FRAME_LEVEL-1:0] fsm_dn_ram_re;
reg [INTER_FRAME_LEVEL-1:0] iter_termination;
reg read_clk, rstn; // shared with all FSMs
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Nets for handshaking protocol between Sys.FSM and Write.FSM
// Input port for Write FSMs from Sys.FSMs
wire [`IB_CNU_DECOMP_funNum-1:0] cnu_wr [0:INTER_FRAME_LEVEL-1];
wire [`IB_VNU_DECOMP_funNum-1:0] vnu_wr [0:INTER_FRAME_LEVEL-1];
wire [INTER_FRAME_LEVEL-1:0] dnu_wr;
// Output port from Write FSMs to Sys.FSMs
wire [`IB_CNU_DECOMP_funNum-1:0] cn_iter_update [0:INTER_FRAME_LEVEL-1];
wire [`IB_VNU_DECOMP_funNum-1:0] vn_iter_update [0:INTER_FRAME_LEVEL-1];
wire [INTER_FRAME_LEVEL-1:0] dn_iter_update;
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Nets of Write.FSMs

wire [2:0] dn_write_fsm_state [0:INTER_FRAME_LEVEL-1];
wire dn_ram_write_en;

// CNU6 Update Iteration Control - Output
wire [`IB_CNU_DECOMP_funNum-1:0] cn_ram_write_en;
wire cn_rom_port_fetch [0:`IB_CNU_DECOMP_funNum-1]; // to enable the ib-map starting to fetch data from read port of IB ROM
wire cn_ram_write_en [0:`IB_CNU_DECOMP_funNum-1];
wire cn_ram_mux_en [0:`IB_CNU_DECOMP_funNum-1];
wire c6ib_rom_rst [0:`IB_CNU_DECOMP_funNum-1];
wire [1:0] cn_write_busy [0:`IB_CNU_DECOMP_funNum-1];
wire [2:0] cn_write_fsm_state [0:INTER_FRAME_LEVEL-1];
// VNU3 Update Iteration Control - Output
wire [`IB_VNU_DECOMP_funNum-1:0] vn_ram_write_en;
wire vn_rom_port_fetch [0:`IB_VNU_DECOMP_funNum-1]; // to enable the ib-map starting to fetch data from read port of IB ROM
wire vn_ram_write_en [0:`IB_VNU_DECOMP_funNum-1];
wire vn_ram_mux_en [0:`IB_VNU_DECOMP_funNum-1];
wire v3ib_rom_rst [0:`IB_VNU_DECOMP_funNum-1];
wire [1:0] vn_write_busy [0:`IB_VNU_DECOMP_funNum-1];
wire [2:0] vn_write_fsm_state [0:INTER_FRAME_LEVEL-1];
// DNU Update Iteration Control - Output
wire dn_ram_write_en;
wire dn_rom_port_fetch; // to enable the ib-map starting to fetch data from read port of IB ROM
wire dn_ram_write_en;
wire dn_ram_mux_en;
wire d3ib_rom_rst;
wire [1:0] dn_write_busy;
wire [2:0] dn_write_fsm_state [0:INTER_FRAME_LEVEL-1];
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Nets of VNU and CNU extrinsic messages
reg [`DATAPATH_WIDTH-1:0] c2v_parallel_in;
reg [`DATAPATH_WIDTH-1:0] v2c_parallel_in;
wire [`DATAPATH_WIDTH-1:0] c2v_parallel_out;
wire [`DATAPATH_WIDTH-1:0] v2c_parallel_out;
wire extrinsic_route; // 1-bit message-passing route
reg c2v_msg_busy; 
reg v2c_msg_busy;
wire c2v_latch_en, v2c_latch_en; 
reg [`DATAPATH_WIDTH-1:0] c2v_latch; // latch the extrinsic message right after PSP which will be fetch by CNU
reg [`DATAPATH_WIDTH-1:0] v2c_latch; // latch the extrinsic message right after PSP which will be fetch by VNU 
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Instantiation of Sys.FSMs
sys_control_unit #(
    //.CNU_PIPELINE_LEVEL  (5-1), // the last pipeline register is actually shared with P2P_C
    //.VNU_PIPELINE_LEVEL  (3-1), // the last pipeline register is actually shared with P2P_V
    .INIT_INTER_FRAME_EN (0)
) frame_fsm_0 (
	// output port for IB-ROM update
	.cnu_wr (cnu_wr[0]),
	.vnu_wr (vnu_wr[0]),
	.dnu_wr (dnu_wr[0]),

    .llr_fetch  (llr_fetch[0]),
    .v2c_src    (v2c_src[0]),
    .v2c_msg_en (v2c_msg_en[0]),
    .cnu_rd     (cnu_rd[0]),
    .c2v_msg_en (c2v_msg_en[0]),
    .vnu_rd     (vnu_rd[0]),
	.dnu_rd		(dnu_rd[0]),
	.c2v_load	(c2v_load[0]), // load enable signal to parallel-to-serial converter
	.v2c_load	(v2c_load[0]), // load enable signal to parallel-to-serial converter
    .inter_frame_en (inter_frame_en[0]),
    .de_frame_start (de_frame_start[0]),
    /*obsoleted*///.cn_ram_re (fsm_cn_ram_re[0]),
    /*obsoleted*///.vn_ram_re (fsm_vn_ram_re[0]),
	/*obsoleted*///.dn_ram_re (fsm_dn_ram_re[0]),
    .state (sys_fsm_state[0]),
    
	// Input port acknowledging from Write/Update FSMs
	.cn_iter_update (cn_iter_update[0]),
	.vn_iter_update (vn_iter_update[0]),
	.dn_iter_update (dn_iter_update[0]),
	
    .termination (iter_termination[0]),
    .inter_frame_align (/*iter_termination[1]*/1'b0),
    .read_clk (read_clk),
    .fsm_en (fsm_en[0]), // enable this FSM only when IB-CNU and VNU RAMs stop write operation
    .rstn (rstn)
);
//and and0(fsm_en[0], rstn, inter_frame_en[1]);

wire decoder_busy;
reg [1:0] next_codeword;
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) fsm_en[0] <= 1'b0;
	else if (codeword_cnt == 0 && iter_cnt == 0) fsm_en[0] <= 1'b1; // to activate in the first time only
	else fsm_en[0] <= ~next_codeword[0];
end
assign decoder_busy = inter_frame_en[0];
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) next_codeword <= 0;
	else next_codeword[1:0] <= {next_codeword[0], iter_termination[0]};
end

/*
sys_control_unit #(
    .CNU_PIPELINE_LEVEL  (5-1), // the last pipeline register is actually shared with P2P_C
    .VNU_PIPELINE_LEVEL  (3-1), // the last pipeline register is actually shared with P2P_V
    .INIT_INTER_FRAME_EN (1)
) frame_fsm_1 (
    .llr_fetch  (llr_fetch[1]),
    .v2c_src    (v2c_src[1]),
    .v2c_msg_en (v2c_msg_en[1]),
    .cnu_rd     (cnu_rd[1]),
    .c2v_msg_en (c2v_msg_en[1]),
    .vnu_rd     (vnu_rd[1]),
    .inter_frame_en (inter_frame_en[1]),
    .de_frame_start (de_frame_start[1]),
    .cn_ram_we (fsm_cn_ram_we[1]),
    .vn_ram_we (fsm_vn_ram_we[1]),
    .state (sys_fsm_state[1]),
    
    .termination (iter_termination[1]),
    .inter_frame_align (iter_termination[0]),
    .read_clk (read_clk),
    .fsm_en (fsm_en[1]), // enable this FSM only when IB-CNU and VNU RAMs stop write operation
    .rstn (rstn)
);
and and1(fsm_en[1], rstn, inter_frame_en[0]);
*/
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Instantiation of Memory System
mem_sys mem_u0(
	// Memory System - Ouput
	.cn_iter0_m0_portA_dout(cn_iter0_m0_portA_dout[CN_RD_BW-1:0]),
	.cn_iter0_m0_portB_dout(cn_iter0_m0_portB_dout[CN_RD_BW-1:0]),
	.cn_iter0_m1_portA_dout(cn_iter0_m1_portA_dout[CN_RD_BW-1:0]),
	.cn_iter0_m1_portB_dout(cn_iter0_m1_portB_dout[CN_RD_BW-1:0]),
	.cn_iter0_m2_portA_dout(cn_iter0_m2_portA_dout[CN_RD_BW-1:0]),
	.cn_iter0_m2_portB_dout(cn_iter0_m2_portB_dout[CN_RD_BW-1:0]),
	.cn_iter0_m3_portA_dout(cn_iter0_m3_portA_dout[CN_RD_BW-1:0]),
	.cn_iter0_m3_portB_dout(cn_iter0_m3_portB_dout[CN_RD_BW-1:0]),
	.cn_iter1_m0_portA_dout(cn_iter1_m0_portA_dout[CN_RD_BW-1:0]),
	.cn_iter1_m0_portB_dout(cn_iter1_m0_portB_dout[CN_RD_BW-1:0]),
	.cn_iter1_m1_portA_dout(cn_iter1_m1_portA_dout[CN_RD_BW-1:0]),
	.cn_iter1_m1_portB_dout(cn_iter1_m1_portB_dout[CN_RD_BW-1:0]),
	.cn_iter1_m2_portA_dout(cn_iter1_m2_portA_dout[CN_RD_BW-1:0]),
	.cn_iter1_m2_portB_dout(cn_iter1_m2_portB_dout[CN_RD_BW-1:0]),
	.cn_iter1_m3_portA_dout(cn_iter1_m3_portA_dout[CN_RD_BW-1:0]),
	.cn_iter1_m3_portB_dout(cn_iter1_m3_portB_dout[CN_RD_BW-1:0]),
	
	.vn_iter0_m0_portA_dout (vn_iter0_m0_portA_dout[VN_RD_BW-1:0]),
	.vn_iter0_m0_portB_dout (vn_iter0_m0_portB_dout[VN_RD_BW-1:0]),
	.vn_iter0_m1_portA_dout (vn_iter0_m1_portA_dout[VN_RD_BW-1:0]),
	.vn_iter0_m1_portB_dout (vn_iter0_m1_portB_dout[VN_RD_BW-1:0]),
	.vn_iter1_m0_portA_dout (vn_iter1_m0_portA_dout[VN_RD_BW-1:0]),
	.vn_iter1_m0_portB_dout (vn_iter1_m0_portB_dout[VN_RD_BW-1:0]),
	.vn_iter1_m1_portA_dout (vn_iter1_m1_portA_dout[VN_RD_BW-1:0]),
	.vn_iter1_m1_portB_dout (vn_iter1_m1_portB_dout[VN_RD_BW-1:0]),
	.dn_iter0_portA_dout (dn_iter0_m2_portA_dout[DN_RD_BW-1:0]),
	.dn_iter0_portB_dout (dn_iter0_m2_portB_dout[DN_RD_BW-1:0]),
	.dn_iter1_portA_dout (dn_iter1_m2_portA_dout[DN_RD_BW-1:0]),
	.dn_iter1_portB_dout (dn_iter1_m2_portB_dout[DN_RD_BW-1:0]),	
	
	// Memory System - Input
	.cn_iter0_m0_portA_addr (cn_rom_read_addrA[0]),
	.cn_iter0_m0_portB_addr (cn_rom_read_addrB[0]),
	.cn_iter0_m1_portA_addr (cn_rom_read_addrA[1]),
	.cn_iter0_m1_portB_addr (cn_rom_read_addrB[1]),
	.cn_iter0_m2_portA_addr (cn_rom_read_addrA[2]),
	.cn_iter0_m2_portB_addr (cn_rom_read_addrB[2]),
	.cn_iter0_m3_portA_addr (cn_rom_read_addrA[3]),
	.cn_iter0_m3_portB_addr (cn_rom_read_addrB[3]),
	.cn_iter1_m0_portA_addr (cn_rom_read_addrA[0]),
	.cn_iter1_m0_portB_addr (cn_rom_read_addrB[0]),
	.cn_iter1_m1_portA_addr (cn_rom_read_addrA[1]),
	.cn_iter1_m1_portB_addr (cn_rom_read_addrB[1]),
	.cn_iter1_m2_portA_addr (cn_rom_read_addrA[2]),
	.cn_iter1_m2_portB_addr (cn_rom_read_addrB[2]),
	.cn_iter1_m3_portA_addr (cn_rom_read_addrA[3]),
	.cn_iter1_m3_portB_addr (cn_rom_read_addrB[3]),
	
	.vn_iter0_m0_portA_addr (vn_rom_read_addrA[0]),
	.vn_iter0_m0_portB_addr (vn_rom_read_addrB[0]),
	.vn_iter0_m1_portA_addr (vn_rom_read_addrA[1]),
	.vn_iter0_m1_portB_addr (vn_rom_read_addrB[1]),
	.vn_iter1_m0_portA_addr (vn_rom_read_addrA[0]),
	.vn_iter1_m0_portB_addr (vn_rom_read_addrB[0]),
	.vn_iter1_m1_portA_addr (vn_rom_read_addrA[1]),
	.vn_iter1_m1_portB_addr (vn_rom_read_addrB[1]),	
	.dn_iter0_portA_addr (dn_rom_read_addrA[ROM_ADDR_BW-1:0]),
	.dn_iter0_portB_addr (dn_rom_read_addrB[ROM_ADDR_BW-1:0]),
	.dn_iter1_portA_addr (dn_rom_read_addrA[ROM_ADDR_BW-1:0]),
	.dn_iter1_portB_addr (dn_rom_read_addrB[ROM_ADDR_BW-1:0]),
	.cn_write_clk (cn_write_clk),
	.vn_write_clk (vn_write_clk),
	.dn_write_clk (dn_write_clk)
);

c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mA0(
	.dout (cn_portA_dout[0]),
	.iter0_din (cn_iter0_m0_portA_dout),
	.iter1_din (cn_iter1_m0_portA_dout),
	.iter_switch (cn_iter_switch[0])
);
c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mA1(
	.dout (cn_portA_dout[1]),
	.iter0_din  (cn_iter0_m1_portA_dout),
	.iter1_din  (cn_iter1_m1_portA_dout),
	.iter_switch (cn_iter_switch[1]) 
);
c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mA2(
	.dout (cn_portA_dout[2]),
	.iter0_din  (cn_iter0_m2_portA_dout),
	.iter1_din  (cn_iter1_m2_portA_dout),
	.iter_switch (cn_iter_switch[2]) 
);
c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mA3(
	.dout (cn_portA_dout[3]),
	.iter0_din  (cn_iter0_m3_portA_dout),
	.iter1_din  (cn_iter1_m3_portA_dout),
	.iter_switch (cn_iter_switch[3]) 
);
c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mB0(
	.dout (cn_portB_dout[0]),
	.iter0_din (cn_iter0_m0_portB_dout),
	.iter1_din (cn_iter1_m0_portB_dout),
	.iter_switch (cn_iter_switch[0])
);
c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mB1(
	.dout (cn_portB_dout[1]),
	.iter0_din  (cn_iter0_m1_portB_dout),
	.iter1_din  (cn_iter1_m1_portB_dout),
	.iter_switch (cn_iter_switch[1]) 
);
c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mB2(
	.dout (cn_portB_dout[2]),
	.iter0_din  (cn_iter0_m2_portB_dout),
	.iter1_din  (cn_iter1_m2_portB_dout),
	.iter_switch (cn_iter_switch[2]) 
);
c6rom_iter_mux #(.ROM_RD_BW(CN_RD_BW)) c6rom_iter_mux_mB3(
	.dout (cn_portB_dout[3]),
	.iter0_din  (cn_iter0_m3_portB_dout),
	.iter1_din  (cn_iter1_m3_portB_dout),
	.iter_switch (cn_iter_switch[3]) 
);

v3rom_iter_mux #(.ROM_RD_BW(VN_RD_BW)) v3rom_iter_mux_mA0(
	.dout        (vn_portA_dout[0]),
	.iter0_din   (vn_iter0_m0_portA_dout),
	.iter1_din   (vn_iter1_m0_portA_dout),
	.iter_switch (vn_iter_switch[0])
);
v3rom_iter_mux #(.ROM_RD_BW(VN_RD_BW)) v3rom_iter_mux_mA1(
	.dout        (vn_portA_dout[1]),
	.iter0_din   (vn_iter0_m1_portA_dout),
	.iter1_din   (vn_iter1_m1_portA_dout),
	.iter_switch (vn_iter_switch[1]) 
);
d3rom_iter_mux #(.ROM_RD_BW(DN_RD_BW)) d3rom_iter_mux_mA2(
	.dout        (dn_portA_dout[DN_RD_BW-1:0]),
	.iter0_din   (dn_iter0_m2_portA_dout[DN_RD_BW-1:0]),
	.iter1_din   (dn_iter1_m2_portA_dout[DN_RD_BW-1:0]),
	.iter_switch (dn_iter_switch) 
);
v3rom_iter_mux #(.ROM_RD_BW(VN_RD_BW)) v3rom_iter_mux_mB0(
	.dout        (vn_portB_dout[0]),
	.iter0_din   (vn_iter0_m0_portB_dout),
	.iter1_din   (vn_iter1_m0_portB_dout),
	.iter_switch (vn_iter_switch[0])
);
v3rom_iter_mux #(.ROM_RD_BW(VN_RD_BW)) v3rom_iter_mux_mB1(
	.dout        (vn_portB_dout[1]),
	.iter0_din   (vn_iter0_m1_portB_dout),
	.iter1_din   (vn_iter1_m1_portB_dout),
	.iter_switch (vn_iter_switch[1]) 
);
d3rom_iter_mux #(.ROM_RD_BW(DN_RD_BW)) d3rom_iter_mux_mB2(
	.dout        (dn_portB_dout[DN_RD_BW-1:0]),
	.iter0_din   (dn_iter0_m2_portB_dout[DN_RD_BW-1:0]),
	.iter1_din   (dn_iter1_m2_portB_dout[DN_RD_BW-1:0]),
	.iter_switch (dn_iter_switch) 
);
//////////////////////////////////////////////////////////////////////////////////////////////////////
// Instantiation of Write.FSMs (for simulation only)
generate
		genvar i, j;
		// For CNUs
		for(i=0;i<`IB_CNU_DECOMP_funNum;i=i+1) begin : cn_wr_fsm_inst		
			cnu6_wr_fsm #(.LOAD_CYCLE(CN_LOAD_CYCLE)) cnu6_wr_fsm_u0 (
				// FSM - Output
				.rom_port_fetch (cn_rom_port_fetch[i]), // to enable the ib-map starting to fetch data from read port of IB ROM
				.ram_write_en   (cn_ram_write_en[i]),
				.ram_mux_en     (cn_ram_mux_en[i]),
				.iter_update    (cn_iter_update[0][i]),
				.c6ib_rom_rst   (c6ib_rom_rst[i]),
				.busy           (cn_write_busy[i]),
				//.state          (cn_write_fsm_state[0]),
				
				// FSM - Input
				.write_clk (cn_write_clk),
				.rstn (/*rstn*/fsm_en[0]),
				.iter_rqst (cnu_wr[0][i]),
				.iter_termination (iter_termination[0])
				//.pipeline_en (pipeline_en[i])	// deprecated
			);
		
			rom_iter_selector #(.ITER_ADDR_BW(ITER_ADDR_BW)) rom_iter_selector_m03(
				.iter_switch (cn_iter_switch[i]),
				.rom_read_addr (cn_rom_read_addrA[i][CN_ROM_ADDR_BW-1:CN_ITER_ADDR_BW]),
				.write_clk (write_clk),
				.rstn (rstn_cnu_fsm[i])
			);
			
			//initial cn_iter_switch[i] <= 1'b0;
			//always @(posedge write_clk) begin
			//	if((rom_read_addrA[i][ROM_ADDR_BW-1:ITER_ADDR_BW] == 5'd24))
			//		cn_iter_switch[i] <= ~cn_iter_switch[i];
			//end
			
			cn_mem_latch #(
				.ROM_RD_BW    (CN_ROM_RD_BW), 
				.ROM_ADDR_BW  (CN_ROM_ADDR_BW),    			    
				.PAGE_ADDR_BW (CN_PAGE_ADDR_BW), 								
				.ITER_ADDR_BW (CN_ITER_ADDR_BW)
			) cn_mem_latch_m03(
				// Memory Latch - Output	
				.latch_outA (cn_latch_outA[i]),
				.latch_outB (cn_latch_outB[i]),
				.rom_read_addrA (cn_rom_read_addrA[i]),
				.rom_read_addrB (cn_rom_read_addrB[i]),
				// Memory Latch - Input 
				.latch_inA (cn_portA_dout[i]),
				.latch_inB (cn_portB_dout[i]),
				.latch_iterA (5'd0), // base address for latch A to indicate the iteration index
				.latch_iterB (5'd0), // base address for latch B to indicate the iteration index
				.rstn (cn_rom_port_fetch[i]), // asserted/deasserted by "rom_port_fetch" signal of Iteration Update Control Unit
				.write_clk (write_clk)
			);
			
			cn_Waddr_counter #(.PAGE_ADDR_BW (CN_PAGE_ADDR_BW)) cn_page_addr_cntM03 (
				.wr_page_addr (cn_wr_page_addr[i]),
				
				.en (cn_ram_write_en[i]),
				.write_clk (write_clk),
				.rstn (~c6ib_rom_rst[i])
			);
		end
		/*----------------------------------------------------------*/
		// For VNUs
		for(j=0;j<`IB_VNU_DECOMP_funNum;j=j+1) begin : vn_wr_fsm_inst
			vnu3_wr_fsm #(.LOAD_CYCLE(VN_LOAD_CYCLE)) vnu3_wr_fsm_u0 (
				// FSM - Output
				.rom_port_fetch (vn_rom_port_fetch[j]), // to enable the ib-map starting to fetch data from read port of IB ROM
				.ram_write_en   (vn_ram_write_en[j]),
				.ram_mux_en     (vn_ram_mux_en[j]),
				.iter_update    (vn_iter_update[0][j]),
				.v3ib_rom_rst   (v3ib_rom_rst[j]),
				.busy           (vn_write_busy[j]),
				//.state (vn_write_fsm_state[0]),
				
				// FSM - Input
				.write_clk (vn_write_clk),
				.rstn (/*rstn*/fsm_en[0]),
				.iter_rqst (vnu_wr[0][j]),
				.iter_termination (iter_termination[0])
				//.pipeline_en (pipeline_en[j])	// deprecated
			);
			v3rom_iter_selector #(.ITER_ADDR_BW(VN_ITER_ADDR_BW)) v3rom_iter_selector_m01(
				.iter_switch   (vn_iter_switch[j]),
				.rom_read_addr (vn_rom_read_addrA[j][VN_ROM_ADDR_BW-1:VN_ITER_ADDR_BW]),
				.write_clk     (write_clk),
				.rstn          (rstn_vnu_fsm[j])
			);
		
			//initial vn_iter_switch[i] <= 1'b0;
			//always @(posedge write_clk) begin
			//	if((vn_rom_read_addrA[i][ROM_ADDR_BW-1:ITER_ADDR_BW] == 5'd24))
			//		vn_iter_switch[i] <= ~vn_iter_switch[i];
			//end
			
			vn_mem_latch #(
				.ROM_RD_BW    (VN_ROM_RD_BW), 
				.ROM_ADDR_BW  (VN_ROM_ADDR_BW),    			    
				.PAGE_ADDR_BW (VN_PAGE_ADDR_BW), 								
				.ITER_ADDR_BW (VN_ITER_ADDR_BW)
			) vn_mem_latch_m01(
				// Memory Latch - Output	
				.latch_outA (vn_latch_outA[j]),
				.latch_outB (vn_latch_outB[j]),
				.rom_read_addrA (vn_rom_read_addrA[j]),
				.rom_read_addrB (vn_rom_read_addrB[j]),
				// Memory Latch - Input 
				.latch_inA (vn_portA_dout[j]),
				.latch_inB (vn_portB_dout[j]),
				.latch_iterA (5'd0), // base address for latch A to indicate the iteration index
				.latch_iterB (5'd0), // base address for latch B to indicate the iteration index
				.rstn (vn_rom_port_fetch[j]), // asserted/deasserted by "rom_port_fetch" signal of Iteration Update Control Unit
				.write_clk (write_clk)
			);

			vn_Waddr_counter #(.PAGE_ADDR_BW (VN_PAGE_ADDR_BW)) vn_page_addr_vntM01 (
				.wr_page_addr (vn_wr_page_addr[j]),
				
				.en (vn_ram_write_en[j]),
				.write_clk (write_clk),
				.rstn (~v3ib_rom_rst[j])
			);
		end
endgenerate
dnu3_wr_fsm #(.LOAD_CYCLE(DN_LOAD_CYCLE)) dnu3_wr_fsm_u0 (
	// FSM - Output
	.rom_port_fetch (dn_rom_port_fetch), // to enable the ib-map starting to fetch data from read port of IB ROM
	.ram_write_en   (dn_ram_write_en),
	.ram_mux_en     (dn_ram_mux_en),
	.iter_update    (dn_iter_update[0]),
	.v3ib_rom_rst   (d3ib_rom_rst),
	.busy           (dn_busy),
	//.state          (dn_write_fsm_state[0]),
	// FSM - Input
	.write_clk        (dn_write_clk),
	.rstn             (/*rstn*/fsm_en[0]),
	.iter_rqst        (dnu_wr[0]),
	.iter_termination (iter_termination[0])
	//.pipeline_en    (vn_pipeline_en[i])	// deprecated
);
dn_mem_latch #(
	.ROM_RD_BW    (DN_ROM_RD_BW), 
	.ROM_ADDR_BW  (DN_ROM_ADDR_BW),    			    
	.PAGE_ADDR_BW (DN_PAGE_ADDR_BW), 								
	.ITER_ADDR_BW (DN_ITER_ADDR_BW)
) dn_mem_latch_m2(
	// Memory Latch - Output	
	.latch_outA (dn_latch_outA[DN_ROM_RD_BW-1:0]),
	.latch_outB (dn_latch_outB[DN_ROM_RD_BW-1:0]),
	.rom_read_addrA (dn_rom_read_addrA[DN_ROM_ADDR_BW-1:0]),
	.rom_read_addrB (dn_rom_read_addrB[DN_ROM_ADDR_BW-1:0]),
	// Memory Latch - Input 
	.latch_inA (dn_portA_dout[DN_RD_BW-1:0]),
	.latch_inB (dn_portB_dout[DN_RD_BW-1:0]),
	.latch_iterA (5'd0), // base address for latch A to indicate the iteration index
	.latch_iterB (5'd0), // base address for latch B to indicate the iteration index
	.rstn (dn_rom_port_fetch), // asserted/deasserted by "rom_port_fetch" signal of Iteration Update Control Unit
	.write_clk (write_clk)
);

dn_Waddr_counter #(.PAGE_ADDR_BW (DN_PAGE_ADDR_BW)) dn_page_addr_vntM2 (
	.wr_page_addr (dn_wr_page_addr[DN_PAGE_ADDR_BW-1:0]),
	
	.en (dn_ram_write_en),
	.write_clk (write_clk),
	.rstn (~d3ib_rom_rst)
);
/*---------------------------------------------------------------------*/
// Instantiation of Routing Network with PSP converter
fully_parallel_route routing_network(
	// (N-K) number of check-to-Variable message buses, each of which is d_c bit width as input ports of this routing network
	.v2c_parallelOut_00(v2c_out0[0]),
	.v2c_parallelOut_01(v2c_out1[0]),
	.v2c_parallelOut_02(v2c_out2[0]),
	.v2c_parallelOut_03(v2c_out3[0]),
	.v2c_parallelOut_04(v2c_out4[0]),
	.v2c_parallelOut_05(v2c_out5[0]),
	.v2c_parallelOut_10(v2c_out0[1]),
	.v2c_parallelOut_11(v2c_out1[1]),
	.v2c_parallelOut_12(v2c_out2[1]),
	.v2c_parallelOut_13(v2c_out3[1]),
	.v2c_parallelOut_14(v2c_out4[1]),
	.v2c_parallelOut_15(v2c_out5[1]),
	.v2c_parallelOut_20(v2c_out0[2]),
	.v2c_parallelOut_21(v2c_out1[2]),
	.v2c_parallelOut_22(v2c_out2[2]),
	.v2c_parallelOut_23(v2c_out3[2]),
	.v2c_parallelOut_24(v2c_out4[2]),
	.v2c_parallelOut_25(v2c_out5[2]),
	.v2c_parallelOut_30(v2c_out0[3]),
	.v2c_parallelOut_31(v2c_out1[3]),
	.v2c_parallelOut_32(v2c_out2[3]),
	.v2c_parallelOut_33(v2c_out3[3]),
	.v2c_parallelOut_34(v2c_out4[3]),
	.v2c_parallelOut_35(v2c_out5[3]),
	.v2c_parallelOut_40(v2c_out0[4]),
	.v2c_parallelOut_41(v2c_out1[4]),
	.v2c_parallelOut_42(v2c_out2[4]),
	.v2c_parallelOut_43(v2c_out3[4]),
	.v2c_parallelOut_44(v2c_out4[4]),
	.v2c_parallelOut_45(v2c_out5[4]),
	.v2c_parallelOut_50(v2c_out0[5]),
	.v2c_parallelOut_51(v2c_out1[5]),
	.v2c_parallelOut_52(v2c_out2[5]),
	.v2c_parallelOut_53(v2c_out3[5]),
	.v2c_parallelOut_54(v2c_out4[5]),
	.v2c_parallelOut_55(v2c_out5[5]),
	.v2c_parallelOut_60(v2c_out0[6]),
	.v2c_parallelOut_61(v2c_out1[6]),
	.v2c_parallelOut_62(v2c_out2[6]),
	.v2c_parallelOut_63(v2c_out3[6]),
	.v2c_parallelOut_64(v2c_out4[6]),
	.v2c_parallelOut_65(v2c_out5[6]),
	.v2c_parallelOut_70(v2c_out0[7]),
	.v2c_parallelOut_71(v2c_out1[7]),
	.v2c_parallelOut_72(v2c_out2[7]),
	.v2c_parallelOut_73(v2c_out3[7]),
	.v2c_parallelOut_74(v2c_out4[7]),
	.v2c_parallelOut_75(v2c_out5[7]),
	.v2c_parallelOut_80(v2c_out0[8]),
	.v2c_parallelOut_81(v2c_out1[8]),
	.v2c_parallelOut_82(v2c_out2[8]),
	.v2c_parallelOut_83(v2c_out3[8]),
	.v2c_parallelOut_84(v2c_out4[8]),
	.v2c_parallelOut_85(v2c_out5[8]),
	.v2c_parallelOut_90(v2c_out0[9]),
	.v2c_parallelOut_91(v2c_out1[9]),
	.v2c_parallelOut_92(v2c_out2[9]),
	.v2c_parallelOut_93(v2c_out3[9]),
	.v2c_parallelOut_94(v2c_out4[9]),
	.v2c_parallelOut_95(v2c_out5[9]),
	.v2c_parallelOut_100(v2c_out0[10]),
	.v2c_parallelOut_101(v2c_out1[10]),
	.v2c_parallelOut_102(v2c_out2[10]),
	.v2c_parallelOut_103(v2c_out3[10]),
	.v2c_parallelOut_104(v2c_out4[10]),
	.v2c_parallelOut_105(v2c_out5[10]),
	.v2c_parallelOut_110(v2c_out0[11]),
	.v2c_parallelOut_111(v2c_out1[11]),
	.v2c_parallelOut_112(v2c_out2[11]),
	.v2c_parallelOut_113(v2c_out3[11]),
	.v2c_parallelOut_114(v2c_out4[11]),
	.v2c_parallelOut_115(v2c_out5[11]),
	.v2c_parallelOut_120(v2c_out0[12]),
	.v2c_parallelOut_121(v2c_out1[12]),
	.v2c_parallelOut_122(v2c_out2[12]),
	.v2c_parallelOut_123(v2c_out3[12]),
	.v2c_parallelOut_124(v2c_out4[12]),
	.v2c_parallelOut_125(v2c_out5[12]),
	.v2c_parallelOut_130(v2c_out0[13]),
	.v2c_parallelOut_131(v2c_out1[13]),
	.v2c_parallelOut_132(v2c_out2[13]),
	.v2c_parallelOut_133(v2c_out3[13]),
	.v2c_parallelOut_134(v2c_out4[13]),
	.v2c_parallelOut_135(v2c_out5[13]),
	.v2c_parallelOut_140(v2c_out0[14]),
	.v2c_parallelOut_141(v2c_out1[14]),
	.v2c_parallelOut_142(v2c_out2[14]),
	.v2c_parallelOut_143(v2c_out3[14]),
	.v2c_parallelOut_144(v2c_out4[14]),
	.v2c_parallelOut_145(v2c_out5[14]),
	.v2c_parallelOut_150(v2c_out0[15]),
	.v2c_parallelOut_151(v2c_out1[15]),
	.v2c_parallelOut_152(v2c_out2[15]),
	.v2c_parallelOut_153(v2c_out3[15]),
	.v2c_parallelOut_154(v2c_out4[15]),
	.v2c_parallelOut_155(v2c_out5[15]),
	.v2c_parallelOut_160(v2c_out0[16]),
	.v2c_parallelOut_161(v2c_out1[16]),
	.v2c_parallelOut_162(v2c_out2[16]),
	.v2c_parallelOut_163(v2c_out3[16]),
	.v2c_parallelOut_164(v2c_out4[16]),
	.v2c_parallelOut_165(v2c_out5[16]),
	.v2c_parallelOut_170(v2c_out0[17]),
	.v2c_parallelOut_171(v2c_out1[17]),
	.v2c_parallelOut_172(v2c_out2[17]),
	.v2c_parallelOut_173(v2c_out3[17]),
	.v2c_parallelOut_174(v2c_out4[17]),
	.v2c_parallelOut_175(v2c_out5[17]),
	.v2c_parallelOut_180(v2c_out0[18]),
	.v2c_parallelOut_181(v2c_out1[18]),
	.v2c_parallelOut_182(v2c_out2[18]),
	.v2c_parallelOut_183(v2c_out3[18]),
	.v2c_parallelOut_184(v2c_out4[18]),
	.v2c_parallelOut_185(v2c_out5[18]),
	.v2c_parallelOut_190(v2c_out0[19]),
	.v2c_parallelOut_191(v2c_out1[19]),
	.v2c_parallelOut_192(v2c_out2[19]),
	.v2c_parallelOut_193(v2c_out3[19]),
	.v2c_parallelOut_194(v2c_out4[19]),
	.v2c_parallelOut_195(v2c_out5[19]),
	.v2c_parallelOut_200(v2c_out0[20]),
	.v2c_parallelOut_201(v2c_out1[20]),
	.v2c_parallelOut_202(v2c_out2[20]),
	.v2c_parallelOut_203(v2c_out3[20]),
	.v2c_parallelOut_204(v2c_out4[20]),
	.v2c_parallelOut_205(v2c_out5[20]),
	.v2c_parallelOut_210(v2c_out0[21]),
	.v2c_parallelOut_211(v2c_out1[21]),
	.v2c_parallelOut_212(v2c_out2[21]),
	.v2c_parallelOut_213(v2c_out3[21]),
	.v2c_parallelOut_214(v2c_out4[21]),
	.v2c_parallelOut_215(v2c_out5[21]),
	.v2c_parallelOut_220(v2c_out0[22]),
	.v2c_parallelOut_221(v2c_out1[22]),
	.v2c_parallelOut_222(v2c_out2[22]),
	.v2c_parallelOut_223(v2c_out3[22]),
	.v2c_parallelOut_224(v2c_out4[22]),
	.v2c_parallelOut_225(v2c_out5[22]),
	.v2c_parallelOut_230(v2c_out0[23]),
	.v2c_parallelOut_231(v2c_out1[23]),
	.v2c_parallelOut_232(v2c_out2[23]),
	.v2c_parallelOut_233(v2c_out3[23]),
	.v2c_parallelOut_234(v2c_out4[23]),
	.v2c_parallelOut_235(v2c_out5[23]),
	.v2c_parallelOut_240(v2c_out0[24]),
	.v2c_parallelOut_241(v2c_out1[24]),
	.v2c_parallelOut_242(v2c_out2[24]),
	.v2c_parallelOut_243(v2c_out3[24]),
	.v2c_parallelOut_244(v2c_out4[24]),
	.v2c_parallelOut_245(v2c_out5[24]),
	.v2c_parallelOut_250(v2c_out0[25]),
	.v2c_parallelOut_251(v2c_out1[25]),
	.v2c_parallelOut_252(v2c_out2[25]),
	.v2c_parallelOut_253(v2c_out3[25]),
	.v2c_parallelOut_254(v2c_out4[25]),
	.v2c_parallelOut_255(v2c_out5[25]),
	.v2c_parallelOut_260(v2c_out0[26]),
	.v2c_parallelOut_261(v2c_out1[26]),
	.v2c_parallelOut_262(v2c_out2[26]),
	.v2c_parallelOut_263(v2c_out3[26]),
	.v2c_parallelOut_264(v2c_out4[26]),
	.v2c_parallelOut_265(v2c_out5[26]),
	.v2c_parallelOut_270(v2c_out0[27]),
	.v2c_parallelOut_271(v2c_out1[27]),
	.v2c_parallelOut_272(v2c_out2[27]),
	.v2c_parallelOut_273(v2c_out3[27]),
	.v2c_parallelOut_274(v2c_out4[27]),
	.v2c_parallelOut_275(v2c_out5[27]),
	.v2c_parallelOut_280(v2c_out0[28]),
	.v2c_parallelOut_281(v2c_out1[28]),
	.v2c_parallelOut_282(v2c_out2[28]),
	.v2c_parallelOut_283(v2c_out3[28]),
	.v2c_parallelOut_284(v2c_out4[28]),
	.v2c_parallelOut_285(v2c_out5[28]),
	.v2c_parallelOut_290(v2c_out0[29]),
	.v2c_parallelOut_291(v2c_out1[29]),
	.v2c_parallelOut_292(v2c_out2[29]),
	.v2c_parallelOut_293(v2c_out3[29]),
	.v2c_parallelOut_294(v2c_out4[29]),
	.v2c_parallelOut_295(v2c_out5[29]),
	.v2c_parallelOut_300(v2c_out0[30]),
	.v2c_parallelOut_301(v2c_out1[30]),
	.v2c_parallelOut_302(v2c_out2[30]),
	.v2c_parallelOut_303(v2c_out3[30]),
	.v2c_parallelOut_304(v2c_out4[30]),
	.v2c_parallelOut_305(v2c_out5[30]),
	.v2c_parallelOut_310(v2c_out0[31]),
	.v2c_parallelOut_311(v2c_out1[31]),
	.v2c_parallelOut_312(v2c_out2[31]),
	.v2c_parallelOut_313(v2c_out3[31]),
	.v2c_parallelOut_314(v2c_out4[31]),
	.v2c_parallelOut_315(v2c_out5[31]),
	.v2c_parallelOut_320(v2c_out0[32]),
	.v2c_parallelOut_321(v2c_out1[32]),
	.v2c_parallelOut_322(v2c_out2[32]),
	.v2c_parallelOut_323(v2c_out3[32]),
	.v2c_parallelOut_324(v2c_out4[32]),
	.v2c_parallelOut_325(v2c_out5[32]),
	.v2c_parallelOut_330(v2c_out0[33]),
	.v2c_parallelOut_331(v2c_out1[33]),
	.v2c_parallelOut_332(v2c_out2[33]),
	.v2c_parallelOut_333(v2c_out3[33]),
	.v2c_parallelOut_334(v2c_out4[33]),
	.v2c_parallelOut_335(v2c_out5[33]),
	.v2c_parallelOut_340(v2c_out0[34]),
	.v2c_parallelOut_341(v2c_out1[34]),
	.v2c_parallelOut_342(v2c_out2[34]),
	.v2c_parallelOut_343(v2c_out3[34]),
	.v2c_parallelOut_344(v2c_out4[34]),
	.v2c_parallelOut_345(v2c_out5[34]),
	.v2c_parallelOut_350(v2c_out0[35]),
	.v2c_parallelOut_351(v2c_out1[35]),
	.v2c_parallelOut_352(v2c_out2[35]),
	.v2c_parallelOut_353(v2c_out3[35]),
	.v2c_parallelOut_354(v2c_out4[35]),
	.v2c_parallelOut_355(v2c_out5[35]),
	.v2c_parallelOut_360(v2c_out0[36]),
	.v2c_parallelOut_361(v2c_out1[36]),
	.v2c_parallelOut_362(v2c_out2[36]),
	.v2c_parallelOut_363(v2c_out3[36]),
	.v2c_parallelOut_364(v2c_out4[36]),
	.v2c_parallelOut_365(v2c_out5[36]),
	.v2c_parallelOut_370(v2c_out0[37]),
	.v2c_parallelOut_371(v2c_out1[37]),
	.v2c_parallelOut_372(v2c_out2[37]),
	.v2c_parallelOut_373(v2c_out3[37]),
	.v2c_parallelOut_374(v2c_out4[37]),
	.v2c_parallelOut_375(v2c_out5[37]),
	.v2c_parallelOut_380(v2c_out0[38]),
	.v2c_parallelOut_381(v2c_out1[38]),
	.v2c_parallelOut_382(v2c_out2[38]),
	.v2c_parallelOut_383(v2c_out3[38]),
	.v2c_parallelOut_384(v2c_out4[38]),
	.v2c_parallelOut_385(v2c_out5[38]),
	.v2c_parallelOut_390(v2c_out0[39]),
	.v2c_parallelOut_391(v2c_out1[39]),
	.v2c_parallelOut_392(v2c_out2[39]),
	.v2c_parallelOut_393(v2c_out3[39]),
	.v2c_parallelOut_394(v2c_out4[39]),
	.v2c_parallelOut_395(v2c_out5[39]),
	.v2c_parallelOut_400(v2c_out0[40]),
	.v2c_parallelOut_401(v2c_out1[40]),
	.v2c_parallelOut_402(v2c_out2[40]),
	.v2c_parallelOut_403(v2c_out3[40]),
	.v2c_parallelOut_404(v2c_out4[40]),
	.v2c_parallelOut_405(v2c_out5[40]),
	.v2c_parallelOut_410(v2c_out0[41]),
	.v2c_parallelOut_411(v2c_out1[41]),
	.v2c_parallelOut_412(v2c_out2[41]),
	.v2c_parallelOut_413(v2c_out3[41]),
	.v2c_parallelOut_414(v2c_out4[41]),
	.v2c_parallelOut_415(v2c_out5[41]),
	.v2c_parallelOut_420(v2c_out0[42]),
	.v2c_parallelOut_421(v2c_out1[42]),
	.v2c_parallelOut_422(v2c_out2[42]),
	.v2c_parallelOut_423(v2c_out3[42]),
	.v2c_parallelOut_424(v2c_out4[42]),
	.v2c_parallelOut_425(v2c_out5[42]),
	.v2c_parallelOut_430(v2c_out0[43]),
	.v2c_parallelOut_431(v2c_out1[43]),
	.v2c_parallelOut_432(v2c_out2[43]),
	.v2c_parallelOut_433(v2c_out3[43]),
	.v2c_parallelOut_434(v2c_out4[43]),
	.v2c_parallelOut_435(v2c_out5[43]),
	.v2c_parallelOut_440(v2c_out0[44]),
	.v2c_parallelOut_441(v2c_out1[44]),
	.v2c_parallelOut_442(v2c_out2[44]),
	.v2c_parallelOut_443(v2c_out3[44]),
	.v2c_parallelOut_444(v2c_out4[44]),
	.v2c_parallelOut_445(v2c_out5[44]),
	.v2c_parallelOut_450(v2c_out0[45]),
	.v2c_parallelOut_451(v2c_out1[45]),
	.v2c_parallelOut_452(v2c_out2[45]),
	.v2c_parallelOut_453(v2c_out3[45]),
	.v2c_parallelOut_454(v2c_out4[45]),
	.v2c_parallelOut_455(v2c_out5[45]),
	.v2c_parallelOut_460(v2c_out0[46]),
	.v2c_parallelOut_461(v2c_out1[46]),
	.v2c_parallelOut_462(v2c_out2[46]),
	.v2c_parallelOut_463(v2c_out3[46]),
	.v2c_parallelOut_464(v2c_out4[46]),
	.v2c_parallelOut_465(v2c_out5[46]),
	.v2c_parallelOut_470(v2c_out0[47]),
	.v2c_parallelOut_471(v2c_out1[47]),
	.v2c_parallelOut_472(v2c_out2[47]),
	.v2c_parallelOut_473(v2c_out3[47]),
	.v2c_parallelOut_474(v2c_out4[47]),
	.v2c_parallelOut_475(v2c_out5[47]),
	.v2c_parallelOut_480(v2c_out0[48]),
	.v2c_parallelOut_481(v2c_out1[48]),
	.v2c_parallelOut_482(v2c_out2[48]),
	.v2c_parallelOut_483(v2c_out3[48]),
	.v2c_parallelOut_484(v2c_out4[48]),
	.v2c_parallelOut_485(v2c_out5[48]),
	.v2c_parallelOut_490(v2c_out0[49]),
	.v2c_parallelOut_491(v2c_out1[49]),
	.v2c_parallelOut_492(v2c_out2[49]),
	.v2c_parallelOut_493(v2c_out3[49]),
	.v2c_parallelOut_494(v2c_out4[49]),
	.v2c_parallelOut_495(v2c_out5[49]),
	.v2c_parallelOut_500(v2c_out0[50]),
	.v2c_parallelOut_501(v2c_out1[50]),
	.v2c_parallelOut_502(v2c_out2[50]),
	.v2c_parallelOut_503(v2c_out3[50]),
	.v2c_parallelOut_504(v2c_out4[50]),
	.v2c_parallelOut_505(v2c_out5[50]),
	.v2c_parallelOut_510(v2c_out0[51]),
	.v2c_parallelOut_511(v2c_out1[51]),
	.v2c_parallelOut_512(v2c_out2[51]),
	.v2c_parallelOut_513(v2c_out3[51]),
	.v2c_parallelOut_514(v2c_out4[51]),
	.v2c_parallelOut_515(v2c_out5[51]),
	.v2c_parallelOut_520(v2c_out0[52]),
	.v2c_parallelOut_521(v2c_out1[52]),
	.v2c_parallelOut_522(v2c_out2[52]),
	.v2c_parallelOut_523(v2c_out3[52]),
	.v2c_parallelOut_524(v2c_out4[52]),
	.v2c_parallelOut_525(v2c_out5[52]),
	.v2c_parallelOut_530(v2c_out0[53]),
	.v2c_parallelOut_531(v2c_out1[53]),
	.v2c_parallelOut_532(v2c_out2[53]),
	.v2c_parallelOut_533(v2c_out3[53]),
	.v2c_parallelOut_534(v2c_out4[53]),
	.v2c_parallelOut_535(v2c_out5[53]),
	.v2c_parallelOut_540(v2c_out0[54]),
	.v2c_parallelOut_541(v2c_out1[54]),
	.v2c_parallelOut_542(v2c_out2[54]),
	.v2c_parallelOut_543(v2c_out3[54]),
	.v2c_parallelOut_544(v2c_out4[54]),
	.v2c_parallelOut_545(v2c_out5[54]),
	.v2c_parallelOut_550(v2c_out0[55]),
	.v2c_parallelOut_551(v2c_out1[55]),
	.v2c_parallelOut_552(v2c_out2[55]),
	.v2c_parallelOut_553(v2c_out3[55]),
	.v2c_parallelOut_554(v2c_out4[55]),
	.v2c_parallelOut_555(v2c_out5[55]),
	.v2c_parallelOut_560(v2c_out0[56]),
	.v2c_parallelOut_561(v2c_out1[56]),
	.v2c_parallelOut_562(v2c_out2[56]),
	.v2c_parallelOut_563(v2c_out3[56]),
	.v2c_parallelOut_564(v2c_out4[56]),
	.v2c_parallelOut_565(v2c_out5[56]),
	.v2c_parallelOut_570(v2c_out0[57]),
	.v2c_parallelOut_571(v2c_out1[57]),
	.v2c_parallelOut_572(v2c_out2[57]),
	.v2c_parallelOut_573(v2c_out3[57]),
	.v2c_parallelOut_574(v2c_out4[57]),
	.v2c_parallelOut_575(v2c_out5[57]),
	.v2c_parallelOut_580(v2c_out0[58]),
	.v2c_parallelOut_581(v2c_out1[58]),
	.v2c_parallelOut_582(v2c_out2[58]),
	.v2c_parallelOut_583(v2c_out3[58]),
	.v2c_parallelOut_584(v2c_out4[58]),
	.v2c_parallelOut_585(v2c_out5[58]),
	.v2c_parallelOut_590(v2c_out0[59]),
	.v2c_parallelOut_591(v2c_out1[59]),
	.v2c_parallelOut_592(v2c_out2[59]),
	.v2c_parallelOut_593(v2c_out3[59]),
	.v2c_parallelOut_594(v2c_out4[59]),
	.v2c_parallelOut_595(v2c_out5[59]),
	.v2c_parallelOut_600(v2c_out0[60]),
	.v2c_parallelOut_601(v2c_out1[60]),
	.v2c_parallelOut_602(v2c_out2[60]),
	.v2c_parallelOut_603(v2c_out3[60]),
	.v2c_parallelOut_604(v2c_out4[60]),
	.v2c_parallelOut_605(v2c_out5[60]),
	.v2c_parallelOut_610(v2c_out0[61]),
	.v2c_parallelOut_611(v2c_out1[61]),
	.v2c_parallelOut_612(v2c_out2[61]),
	.v2c_parallelOut_613(v2c_out3[61]),
	.v2c_parallelOut_614(v2c_out4[61]),
	.v2c_parallelOut_615(v2c_out5[61]),
	.v2c_parallelOut_620(v2c_out0[62]),
	.v2c_parallelOut_621(v2c_out1[62]),
	.v2c_parallelOut_622(v2c_out2[62]),
	.v2c_parallelOut_623(v2c_out3[62]),
	.v2c_parallelOut_624(v2c_out4[62]),
	.v2c_parallelOut_625(v2c_out5[62]),
	.v2c_parallelOut_630(v2c_out0[63]),
	.v2c_parallelOut_631(v2c_out1[63]),
	.v2c_parallelOut_632(v2c_out2[63]),
	.v2c_parallelOut_633(v2c_out3[63]),
	.v2c_parallelOut_634(v2c_out4[63]),
	.v2c_parallelOut_635(v2c_out5[63]),
	.v2c_parallelOut_640(v2c_out0[64]),
	.v2c_parallelOut_641(v2c_out1[64]),
	.v2c_parallelOut_642(v2c_out2[64]),
	.v2c_parallelOut_643(v2c_out3[64]),
	.v2c_parallelOut_644(v2c_out4[64]),
	.v2c_parallelOut_645(v2c_out5[64]),
	.v2c_parallelOut_650(v2c_out0[65]),
	.v2c_parallelOut_651(v2c_out1[65]),
	.v2c_parallelOut_652(v2c_out2[65]),
	.v2c_parallelOut_653(v2c_out3[65]),
	.v2c_parallelOut_654(v2c_out4[65]),
	.v2c_parallelOut_655(v2c_out5[65]),
	.v2c_parallelOut_660(v2c_out0[66]),
	.v2c_parallelOut_661(v2c_out1[66]),
	.v2c_parallelOut_662(v2c_out2[66]),
	.v2c_parallelOut_663(v2c_out3[66]),
	.v2c_parallelOut_664(v2c_out4[66]),
	.v2c_parallelOut_665(v2c_out5[66]),
	.v2c_parallelOut_670(v2c_out0[67]),
	.v2c_parallelOut_671(v2c_out1[67]),
	.v2c_parallelOut_672(v2c_out2[67]),
	.v2c_parallelOut_673(v2c_out3[67]),
	.v2c_parallelOut_674(v2c_out4[67]),
	.v2c_parallelOut_675(v2c_out5[67]),
	.v2c_parallelOut_680(v2c_out0[68]),
	.v2c_parallelOut_681(v2c_out1[68]),
	.v2c_parallelOut_682(v2c_out2[68]),
	.v2c_parallelOut_683(v2c_out3[68]),
	.v2c_parallelOut_684(v2c_out4[68]),
	.v2c_parallelOut_685(v2c_out5[68]),
	.v2c_parallelOut_690(v2c_out0[69]),
	.v2c_parallelOut_691(v2c_out1[69]),
	.v2c_parallelOut_692(v2c_out2[69]),
	.v2c_parallelOut_693(v2c_out3[69]),
	.v2c_parallelOut_694(v2c_out4[69]),
	.v2c_parallelOut_695(v2c_out5[69]),
	.v2c_parallelOut_700(v2c_out0[70]),
	.v2c_parallelOut_701(v2c_out1[70]),
	.v2c_parallelOut_702(v2c_out2[70]),
	.v2c_parallelOut_703(v2c_out3[70]),
	.v2c_parallelOut_704(v2c_out4[70]),
	.v2c_parallelOut_705(v2c_out5[70]),
	.v2c_parallelOut_710(v2c_out0[71]),
	.v2c_parallelOut_711(v2c_out1[71]),
	.v2c_parallelOut_712(v2c_out2[71]),
	.v2c_parallelOut_713(v2c_out3[71]),
	.v2c_parallelOut_714(v2c_out4[71]),
	.v2c_parallelOut_715(v2c_out5[71]),
	.v2c_parallelOut_720(v2c_out0[72]),
	.v2c_parallelOut_721(v2c_out1[72]),
	.v2c_parallelOut_722(v2c_out2[72]),
	.v2c_parallelOut_723(v2c_out3[72]),
	.v2c_parallelOut_724(v2c_out4[72]),
	.v2c_parallelOut_725(v2c_out5[72]),
	.v2c_parallelOut_730(v2c_out0[73]),
	.v2c_parallelOut_731(v2c_out1[73]),
	.v2c_parallelOut_732(v2c_out2[73]),
	.v2c_parallelOut_733(v2c_out3[73]),
	.v2c_parallelOut_734(v2c_out4[73]),
	.v2c_parallelOut_735(v2c_out5[73]),
	.v2c_parallelOut_740(v2c_out0[74]),
	.v2c_parallelOut_741(v2c_out1[74]),
	.v2c_parallelOut_742(v2c_out2[74]),
	.v2c_parallelOut_743(v2c_out3[74]),
	.v2c_parallelOut_744(v2c_out4[74]),
	.v2c_parallelOut_745(v2c_out5[74]),
	.v2c_parallelOut_750(v2c_out0[75]),
	.v2c_parallelOut_751(v2c_out1[75]),
	.v2c_parallelOut_752(v2c_out2[75]),
	.v2c_parallelOut_753(v2c_out3[75]),
	.v2c_parallelOut_754(v2c_out4[75]),
	.v2c_parallelOut_755(v2c_out5[75]),
	.v2c_parallelOut_760(v2c_out0[76]),
	.v2c_parallelOut_761(v2c_out1[76]),
	.v2c_parallelOut_762(v2c_out2[76]),
	.v2c_parallelOut_763(v2c_out3[76]),
	.v2c_parallelOut_764(v2c_out4[76]),
	.v2c_parallelOut_765(v2c_out5[76]),
	.v2c_parallelOut_770(v2c_out0[77]),
	.v2c_parallelOut_771(v2c_out1[77]),
	.v2c_parallelOut_772(v2c_out2[77]),
	.v2c_parallelOut_773(v2c_out3[77]),
	.v2c_parallelOut_774(v2c_out4[77]),
	.v2c_parallelOut_775(v2c_out5[77]),
	.v2c_parallelOut_780(v2c_out0[78]),
	.v2c_parallelOut_781(v2c_out1[78]),
	.v2c_parallelOut_782(v2c_out2[78]),
	.v2c_parallelOut_783(v2c_out3[78]),
	.v2c_parallelOut_784(v2c_out4[78]),
	.v2c_parallelOut_785(v2c_out5[78]),
	.v2c_parallelOut_790(v2c_out0[79]),
	.v2c_parallelOut_791(v2c_out1[79]),
	.v2c_parallelOut_792(v2c_out2[79]),
	.v2c_parallelOut_793(v2c_out3[79]),
	.v2c_parallelOut_794(v2c_out4[79]),
	.v2c_parallelOut_795(v2c_out5[79]),
	.v2c_parallelOut_800(v2c_out0[80]),
	.v2c_parallelOut_801(v2c_out1[80]),
	.v2c_parallelOut_802(v2c_out2[80]),
	.v2c_parallelOut_803(v2c_out3[80]),
	.v2c_parallelOut_804(v2c_out4[80]),
	.v2c_parallelOut_805(v2c_out5[80]),
	.v2c_parallelOut_810(v2c_out0[81]),
	.v2c_parallelOut_811(v2c_out1[81]),
	.v2c_parallelOut_812(v2c_out2[81]),
	.v2c_parallelOut_813(v2c_out3[81]),
	.v2c_parallelOut_814(v2c_out4[81]),
	.v2c_parallelOut_815(v2c_out5[81]),
	.v2c_parallelOut_820(v2c_out0[82]),
	.v2c_parallelOut_821(v2c_out1[82]),
	.v2c_parallelOut_822(v2c_out2[82]),
	.v2c_parallelOut_823(v2c_out3[82]),
	.v2c_parallelOut_824(v2c_out4[82]),
	.v2c_parallelOut_825(v2c_out5[82]),
	.v2c_parallelOut_830(v2c_out0[83]),
	.v2c_parallelOut_831(v2c_out1[83]),
	.v2c_parallelOut_832(v2c_out2[83]),
	.v2c_parallelOut_833(v2c_out3[83]),
	.v2c_parallelOut_834(v2c_out4[83]),
	.v2c_parallelOut_835(v2c_out5[83]),
	.v2c_parallelOut_840(v2c_out0[84]),
	.v2c_parallelOut_841(v2c_out1[84]),
	.v2c_parallelOut_842(v2c_out2[84]),
	.v2c_parallelOut_843(v2c_out3[84]),
	.v2c_parallelOut_844(v2c_out4[84]),
	.v2c_parallelOut_845(v2c_out5[84]),
	.v2c_parallelOut_850(v2c_out0[85]),
	.v2c_parallelOut_851(v2c_out1[85]),
	.v2c_parallelOut_852(v2c_out2[85]),
	.v2c_parallelOut_853(v2c_out3[85]),
	.v2c_parallelOut_854(v2c_out4[85]),
	.v2c_parallelOut_855(v2c_out5[85]),
	.v2c_parallelOut_860(v2c_out0[86]),
	.v2c_parallelOut_861(v2c_out1[86]),
	.v2c_parallelOut_862(v2c_out2[86]),
	.v2c_parallelOut_863(v2c_out3[86]),
	.v2c_parallelOut_864(v2c_out4[86]),
	.v2c_parallelOut_865(v2c_out5[86]),
	.v2c_parallelOut_870(v2c_out0[87]),
	.v2c_parallelOut_871(v2c_out1[87]),
	.v2c_parallelOut_872(v2c_out2[87]),
	.v2c_parallelOut_873(v2c_out3[87]),
	.v2c_parallelOut_874(v2c_out4[87]),
	.v2c_parallelOut_875(v2c_out5[87]),
	.v2c_parallelOut_880(v2c_out0[88]),
	.v2c_parallelOut_881(v2c_out1[88]),
	.v2c_parallelOut_882(v2c_out2[88]),
	.v2c_parallelOut_883(v2c_out3[88]),
	.v2c_parallelOut_884(v2c_out4[88]),
	.v2c_parallelOut_885(v2c_out5[88]),
	.v2c_parallelOut_890(v2c_out0[89]),
	.v2c_parallelOut_891(v2c_out1[89]),
	.v2c_parallelOut_892(v2c_out2[89]),
	.v2c_parallelOut_893(v2c_out3[89]),
	.v2c_parallelOut_894(v2c_out4[89]),
	.v2c_parallelOut_895(v2c_out5[89]),
	.v2c_parallelOut_900(v2c_out0[90]),
	.v2c_parallelOut_901(v2c_out1[90]),
	.v2c_parallelOut_902(v2c_out2[90]),
	.v2c_parallelOut_903(v2c_out3[90]),
	.v2c_parallelOut_904(v2c_out4[90]),
	.v2c_parallelOut_905(v2c_out5[90]),
	.v2c_parallelOut_910(v2c_out0[91]),
	.v2c_parallelOut_911(v2c_out1[91]),
	.v2c_parallelOut_912(v2c_out2[91]),
	.v2c_parallelOut_913(v2c_out3[91]),
	.v2c_parallelOut_914(v2c_out4[91]),
	.v2c_parallelOut_915(v2c_out5[91]),
	.v2c_parallelOut_920(v2c_out0[92]),
	.v2c_parallelOut_921(v2c_out1[92]),
	.v2c_parallelOut_922(v2c_out2[92]),
	.v2c_parallelOut_923(v2c_out3[92]),
	.v2c_parallelOut_924(v2c_out4[92]),
	.v2c_parallelOut_925(v2c_out5[92]),
	.v2c_parallelOut_930(v2c_out0[93]),
	.v2c_parallelOut_931(v2c_out1[93]),
	.v2c_parallelOut_932(v2c_out2[93]),
	.v2c_parallelOut_933(v2c_out3[93]),
	.v2c_parallelOut_934(v2c_out4[93]),
	.v2c_parallelOut_935(v2c_out5[93]),
	.v2c_parallelOut_940(v2c_out0[94]),
	.v2c_parallelOut_941(v2c_out1[94]),
	.v2c_parallelOut_942(v2c_out2[94]),
	.v2c_parallelOut_943(v2c_out3[94]),
	.v2c_parallelOut_944(v2c_out4[94]),
	.v2c_parallelOut_945(v2c_out5[94]),
	.v2c_parallelOut_950(v2c_out0[95]),
	.v2c_parallelOut_951(v2c_out1[95]),
	.v2c_parallelOut_952(v2c_out2[95]),
	.v2c_parallelOut_953(v2c_out3[95]),
	.v2c_parallelOut_954(v2c_out4[95]),
	.v2c_parallelOut_955(v2c_out5[95]),
	.v2c_parallelOut_960(v2c_out0[96]),
	.v2c_parallelOut_961(v2c_out1[96]),
	.v2c_parallelOut_962(v2c_out2[96]),
	.v2c_parallelOut_963(v2c_out3[96]),
	.v2c_parallelOut_964(v2c_out4[96]),
	.v2c_parallelOut_965(v2c_out5[96]),
	.v2c_parallelOut_970(v2c_out0[97]),
	.v2c_parallelOut_971(v2c_out1[97]),
	.v2c_parallelOut_972(v2c_out2[97]),
	.v2c_parallelOut_973(v2c_out3[97]),
	.v2c_parallelOut_974(v2c_out4[97]),
	.v2c_parallelOut_975(v2c_out5[97]),
	.v2c_parallelOut_980(v2c_out0[98]),
	.v2c_parallelOut_981(v2c_out1[98]),
	.v2c_parallelOut_982(v2c_out2[98]),
	.v2c_parallelOut_983(v2c_out3[98]),
	.v2c_parallelOut_984(v2c_out4[98]),
	.v2c_parallelOut_985(v2c_out5[98]),
	.v2c_parallelOut_990(v2c_out0[99]),
	.v2c_parallelOut_991(v2c_out1[99]),
	.v2c_parallelOut_992(v2c_out2[99]),
	.v2c_parallelOut_993(v2c_out3[99]),
	.v2c_parallelOut_994(v2c_out4[99]),
	.v2c_parallelOut_995(v2c_out5[99]),
	.v2c_parallelOut_1000(v2c_out0[100]),
	.v2c_parallelOut_1001(v2c_out1[100]),
	.v2c_parallelOut_1002(v2c_out2[100]),
	.v2c_parallelOut_1003(v2c_out3[100]),
	.v2c_parallelOut_1004(v2c_out4[100]),
	.v2c_parallelOut_1005(v2c_out5[100]),
	.v2c_parallelOut_1010(v2c_out0[101]),
	.v2c_parallelOut_1011(v2c_out1[101]),
	.v2c_parallelOut_1012(v2c_out2[101]),
	.v2c_parallelOut_1013(v2c_out3[101]),
	.v2c_parallelOut_1014(v2c_out4[101]),
	.v2c_parallelOut_1015(v2c_out5[101]),
	
	// N number of check-to-Variable message buses, each of which is d_v bit width outgoing to serial-to-parallel converters
	.c2v_parallelOut_00(c2v_out0[0]),
	.c2v_parallelOut_01(c2v_out1[0]),
	.c2v_parallelOut_02(c2v_out2[0]),
	.c2v_parallelOut_10(c2v_out0[1]),
	.c2v_parallelOut_11(c2v_out1[1]),
	.c2v_parallelOut_12(c2v_out2[1]),
	.c2v_parallelOut_20(c2v_out0[2]),
	.c2v_parallelOut_21(c2v_out1[2]),
	.c2v_parallelOut_22(c2v_out2[2]),
	.c2v_parallelOut_30(c2v_out0[3]),
	.c2v_parallelOut_31(c2v_out1[3]),
	.c2v_parallelOut_32(c2v_out2[3]),
	.c2v_parallelOut_40(c2v_out0[4]),
	.c2v_parallelOut_41(c2v_out1[4]),
	.c2v_parallelOut_42(c2v_out2[4]),
	.c2v_parallelOut_50(c2v_out0[5]),
	.c2v_parallelOut_51(c2v_out1[5]),
	.c2v_parallelOut_52(c2v_out2[5]),
	.c2v_parallelOut_60(c2v_out0[6]),
	.c2v_parallelOut_61(c2v_out1[6]),
	.c2v_parallelOut_62(c2v_out2[6]),
	.c2v_parallelOut_70(c2v_out0[7]),
	.c2v_parallelOut_71(c2v_out1[7]),
	.c2v_parallelOut_72(c2v_out2[7]),
	.c2v_parallelOut_80(c2v_out0[8]),
	.c2v_parallelOut_81(c2v_out1[8]),
	.c2v_parallelOut_82(c2v_out2[8]),
	.c2v_parallelOut_90(c2v_out0[9]),
	.c2v_parallelOut_91(c2v_out1[9]),
	.c2v_parallelOut_92(c2v_out2[9]),
	.c2v_parallelOut_100(c2v_out0[10]),
	.c2v_parallelOut_101(c2v_out1[10]),
	.c2v_parallelOut_102(c2v_out2[10]),
	.c2v_parallelOut_110(c2v_out0[11]),
	.c2v_parallelOut_111(c2v_out1[11]),
	.c2v_parallelOut_112(c2v_out2[11]),
	.c2v_parallelOut_120(c2v_out0[12]),
	.c2v_parallelOut_121(c2v_out1[12]),
	.c2v_parallelOut_122(c2v_out2[12]),
	.c2v_parallelOut_130(c2v_out0[13]),
	.c2v_parallelOut_131(c2v_out1[13]),
	.c2v_parallelOut_132(c2v_out2[13]),
	.c2v_parallelOut_140(c2v_out0[14]),
	.c2v_parallelOut_141(c2v_out1[14]),
	.c2v_parallelOut_142(c2v_out2[14]),
	.c2v_parallelOut_150(c2v_out0[15]),
	.c2v_parallelOut_151(c2v_out1[15]),
	.c2v_parallelOut_152(c2v_out2[15]),
	.c2v_parallelOut_160(c2v_out0[16]),
	.c2v_parallelOut_161(c2v_out1[16]),
	.c2v_parallelOut_162(c2v_out2[16]),
	.c2v_parallelOut_170(c2v_out0[17]),
	.c2v_parallelOut_171(c2v_out1[17]),
	.c2v_parallelOut_172(c2v_out2[17]),
	.c2v_parallelOut_180(c2v_out0[18]),
	.c2v_parallelOut_181(c2v_out1[18]),
	.c2v_parallelOut_182(c2v_out2[18]),
	.c2v_parallelOut_190(c2v_out0[19]),
	.c2v_parallelOut_191(c2v_out1[19]),
	.c2v_parallelOut_192(c2v_out2[19]),
	.c2v_parallelOut_200(c2v_out0[20]),
	.c2v_parallelOut_201(c2v_out1[20]),
	.c2v_parallelOut_202(c2v_out2[20]),
	.c2v_parallelOut_210(c2v_out0[21]),
	.c2v_parallelOut_211(c2v_out1[21]),
	.c2v_parallelOut_212(c2v_out2[21]),
	.c2v_parallelOut_220(c2v_out0[22]),
	.c2v_parallelOut_221(c2v_out1[22]),
	.c2v_parallelOut_222(c2v_out2[22]),
	.c2v_parallelOut_230(c2v_out0[23]),
	.c2v_parallelOut_231(c2v_out1[23]),
	.c2v_parallelOut_232(c2v_out2[23]),
	.c2v_parallelOut_240(c2v_out0[24]),
	.c2v_parallelOut_241(c2v_out1[24]),
	.c2v_parallelOut_242(c2v_out2[24]),
	.c2v_parallelOut_250(c2v_out0[25]),
	.c2v_parallelOut_251(c2v_out1[25]),
	.c2v_parallelOut_252(c2v_out2[25]),
	.c2v_parallelOut_260(c2v_out0[26]),
	.c2v_parallelOut_261(c2v_out1[26]),
	.c2v_parallelOut_262(c2v_out2[26]),
	.c2v_parallelOut_270(c2v_out0[27]),
	.c2v_parallelOut_271(c2v_out1[27]),
	.c2v_parallelOut_272(c2v_out2[27]),
	.c2v_parallelOut_280(c2v_out0[28]),
	.c2v_parallelOut_281(c2v_out1[28]),
	.c2v_parallelOut_282(c2v_out2[28]),
	.c2v_parallelOut_290(c2v_out0[29]),
	.c2v_parallelOut_291(c2v_out1[29]),
	.c2v_parallelOut_292(c2v_out2[29]),
	.c2v_parallelOut_300(c2v_out0[30]),
	.c2v_parallelOut_301(c2v_out1[30]),
	.c2v_parallelOut_302(c2v_out2[30]),
	.c2v_parallelOut_310(c2v_out0[31]),
	.c2v_parallelOut_311(c2v_out1[31]),
	.c2v_parallelOut_312(c2v_out2[31]),
	.c2v_parallelOut_320(c2v_out0[32]),
	.c2v_parallelOut_321(c2v_out1[32]),
	.c2v_parallelOut_322(c2v_out2[32]),
	.c2v_parallelOut_330(c2v_out0[33]),
	.c2v_parallelOut_331(c2v_out1[33]),
	.c2v_parallelOut_332(c2v_out2[33]),
	.c2v_parallelOut_340(c2v_out0[34]),
	.c2v_parallelOut_341(c2v_out1[34]),
	.c2v_parallelOut_342(c2v_out2[34]),
	.c2v_parallelOut_350(c2v_out0[35]),
	.c2v_parallelOut_351(c2v_out1[35]),
	.c2v_parallelOut_352(c2v_out2[35]),
	.c2v_parallelOut_360(c2v_out0[36]),
	.c2v_parallelOut_361(c2v_out1[36]),
	.c2v_parallelOut_362(c2v_out2[36]),
	.c2v_parallelOut_370(c2v_out0[37]),
	.c2v_parallelOut_371(c2v_out1[37]),
	.c2v_parallelOut_372(c2v_out2[37]),
	.c2v_parallelOut_380(c2v_out0[38]),
	.c2v_parallelOut_381(c2v_out1[38]),
	.c2v_parallelOut_382(c2v_out2[38]),
	.c2v_parallelOut_390(c2v_out0[39]),
	.c2v_parallelOut_391(c2v_out1[39]),
	.c2v_parallelOut_392(c2v_out2[39]),
	.c2v_parallelOut_400(c2v_out0[40]),
	.c2v_parallelOut_401(c2v_out1[40]),
	.c2v_parallelOut_402(c2v_out2[40]),
	.c2v_parallelOut_410(c2v_out0[41]),
	.c2v_parallelOut_411(c2v_out1[41]),
	.c2v_parallelOut_412(c2v_out2[41]),
	.c2v_parallelOut_420(c2v_out0[42]),
	.c2v_parallelOut_421(c2v_out1[42]),
	.c2v_parallelOut_422(c2v_out2[42]),
	.c2v_parallelOut_430(c2v_out0[43]),
	.c2v_parallelOut_431(c2v_out1[43]),
	.c2v_parallelOut_432(c2v_out2[43]),
	.c2v_parallelOut_440(c2v_out0[44]),
	.c2v_parallelOut_441(c2v_out1[44]),
	.c2v_parallelOut_442(c2v_out2[44]),
	.c2v_parallelOut_450(c2v_out0[45]),
	.c2v_parallelOut_451(c2v_out1[45]),
	.c2v_parallelOut_452(c2v_out2[45]),
	.c2v_parallelOut_460(c2v_out0[46]),
	.c2v_parallelOut_461(c2v_out1[46]),
	.c2v_parallelOut_462(c2v_out2[46]),
	.c2v_parallelOut_470(c2v_out0[47]),
	.c2v_parallelOut_471(c2v_out1[47]),
	.c2v_parallelOut_472(c2v_out2[47]),
	.c2v_parallelOut_480(c2v_out0[48]),
	.c2v_parallelOut_481(c2v_out1[48]),
	.c2v_parallelOut_482(c2v_out2[48]),
	.c2v_parallelOut_490(c2v_out0[49]),
	.c2v_parallelOut_491(c2v_out1[49]),
	.c2v_parallelOut_492(c2v_out2[49]),
	.c2v_parallelOut_500(c2v_out0[50]),
	.c2v_parallelOut_501(c2v_out1[50]),
	.c2v_parallelOut_502(c2v_out2[50]),
	.c2v_parallelOut_510(c2v_out0[51]),
	.c2v_parallelOut_511(c2v_out1[51]),
	.c2v_parallelOut_512(c2v_out2[51]),
	.c2v_parallelOut_520(c2v_out0[52]),
	.c2v_parallelOut_521(c2v_out1[52]),
	.c2v_parallelOut_522(c2v_out2[52]),
	.c2v_parallelOut_530(c2v_out0[53]),
	.c2v_parallelOut_531(c2v_out1[53]),
	.c2v_parallelOut_532(c2v_out2[53]),
	.c2v_parallelOut_540(c2v_out0[54]),
	.c2v_parallelOut_541(c2v_out1[54]),
	.c2v_parallelOut_542(c2v_out2[54]),
	.c2v_parallelOut_550(c2v_out0[55]),
	.c2v_parallelOut_551(c2v_out1[55]),
	.c2v_parallelOut_552(c2v_out2[55]),
	.c2v_parallelOut_560(c2v_out0[56]),
	.c2v_parallelOut_561(c2v_out1[56]),
	.c2v_parallelOut_562(c2v_out2[56]),
	.c2v_parallelOut_570(c2v_out0[57]),
	.c2v_parallelOut_571(c2v_out1[57]),
	.c2v_parallelOut_572(c2v_out2[57]),
	.c2v_parallelOut_580(c2v_out0[58]),
	.c2v_parallelOut_581(c2v_out1[58]),
	.c2v_parallelOut_582(c2v_out2[58]),
	.c2v_parallelOut_590(c2v_out0[59]),
	.c2v_parallelOut_591(c2v_out1[59]),
	.c2v_parallelOut_592(c2v_out2[59]),
	.c2v_parallelOut_600(c2v_out0[60]),
	.c2v_parallelOut_601(c2v_out1[60]),
	.c2v_parallelOut_602(c2v_out2[60]),
	.c2v_parallelOut_610(c2v_out0[61]),
	.c2v_parallelOut_611(c2v_out1[61]),
	.c2v_parallelOut_612(c2v_out2[61]),
	.c2v_parallelOut_620(c2v_out0[62]),
	.c2v_parallelOut_621(c2v_out1[62]),
	.c2v_parallelOut_622(c2v_out2[62]),
	.c2v_parallelOut_630(c2v_out0[63]),
	.c2v_parallelOut_631(c2v_out1[63]),
	.c2v_parallelOut_632(c2v_out2[63]),
	.c2v_parallelOut_640(c2v_out0[64]),
	.c2v_parallelOut_641(c2v_out1[64]),
	.c2v_parallelOut_642(c2v_out2[64]),
	.c2v_parallelOut_650(c2v_out0[65]),
	.c2v_parallelOut_651(c2v_out1[65]),
	.c2v_parallelOut_652(c2v_out2[65]),
	.c2v_parallelOut_660(c2v_out0[66]),
	.c2v_parallelOut_661(c2v_out1[66]),
	.c2v_parallelOut_662(c2v_out2[66]),
	.c2v_parallelOut_670(c2v_out0[67]),
	.c2v_parallelOut_671(c2v_out1[67]),
	.c2v_parallelOut_672(c2v_out2[67]),
	.c2v_parallelOut_680(c2v_out0[68]),
	.c2v_parallelOut_681(c2v_out1[68]),
	.c2v_parallelOut_682(c2v_out2[68]),
	.c2v_parallelOut_690(c2v_out0[69]),
	.c2v_parallelOut_691(c2v_out1[69]),
	.c2v_parallelOut_692(c2v_out2[69]),
	.c2v_parallelOut_700(c2v_out0[70]),
	.c2v_parallelOut_701(c2v_out1[70]),
	.c2v_parallelOut_702(c2v_out2[70]),
	.c2v_parallelOut_710(c2v_out0[71]),
	.c2v_parallelOut_711(c2v_out1[71]),
	.c2v_parallelOut_712(c2v_out2[71]),
	.c2v_parallelOut_720(c2v_out0[72]),
	.c2v_parallelOut_721(c2v_out1[72]),
	.c2v_parallelOut_722(c2v_out2[72]),
	.c2v_parallelOut_730(c2v_out0[73]),
	.c2v_parallelOut_731(c2v_out1[73]),
	.c2v_parallelOut_732(c2v_out2[73]),
	.c2v_parallelOut_740(c2v_out0[74]),
	.c2v_parallelOut_741(c2v_out1[74]),
	.c2v_parallelOut_742(c2v_out2[74]),
	.c2v_parallelOut_750(c2v_out0[75]),
	.c2v_parallelOut_751(c2v_out1[75]),
	.c2v_parallelOut_752(c2v_out2[75]),
	.c2v_parallelOut_760(c2v_out0[76]),
	.c2v_parallelOut_761(c2v_out1[76]),
	.c2v_parallelOut_762(c2v_out2[76]),
	.c2v_parallelOut_770(c2v_out0[77]),
	.c2v_parallelOut_771(c2v_out1[77]),
	.c2v_parallelOut_772(c2v_out2[77]),
	.c2v_parallelOut_780(c2v_out0[78]),
	.c2v_parallelOut_781(c2v_out1[78]),
	.c2v_parallelOut_782(c2v_out2[78]),
	.c2v_parallelOut_790(c2v_out0[79]),
	.c2v_parallelOut_791(c2v_out1[79]),
	.c2v_parallelOut_792(c2v_out2[79]),
	.c2v_parallelOut_800(c2v_out0[80]),
	.c2v_parallelOut_801(c2v_out1[80]),
	.c2v_parallelOut_802(c2v_out2[80]),
	.c2v_parallelOut_810(c2v_out0[81]),
	.c2v_parallelOut_811(c2v_out1[81]),
	.c2v_parallelOut_812(c2v_out2[81]),
	.c2v_parallelOut_820(c2v_out0[82]),
	.c2v_parallelOut_821(c2v_out1[82]),
	.c2v_parallelOut_822(c2v_out2[82]),
	.c2v_parallelOut_830(c2v_out0[83]),
	.c2v_parallelOut_831(c2v_out1[83]),
	.c2v_parallelOut_832(c2v_out2[83]),
	.c2v_parallelOut_840(c2v_out0[84]),
	.c2v_parallelOut_841(c2v_out1[84]),
	.c2v_parallelOut_842(c2v_out2[84]),
	.c2v_parallelOut_850(c2v_out0[85]),
	.c2v_parallelOut_851(c2v_out1[85]),
	.c2v_parallelOut_852(c2v_out2[85]),
	.c2v_parallelOut_860(c2v_out0[86]),
	.c2v_parallelOut_861(c2v_out1[86]),
	.c2v_parallelOut_862(c2v_out2[86]),
	.c2v_parallelOut_870(c2v_out0[87]),
	.c2v_parallelOut_871(c2v_out1[87]),
	.c2v_parallelOut_872(c2v_out2[87]),
	.c2v_parallelOut_880(c2v_out0[88]),
	.c2v_parallelOut_881(c2v_out1[88]),
	.c2v_parallelOut_882(c2v_out2[88]),
	.c2v_parallelOut_890(c2v_out0[89]),
	.c2v_parallelOut_891(c2v_out1[89]),
	.c2v_parallelOut_892(c2v_out2[89]),
	.c2v_parallelOut_900(c2v_out0[90]),
	.c2v_parallelOut_901(c2v_out1[90]),
	.c2v_parallelOut_902(c2v_out2[90]),
	.c2v_parallelOut_910(c2v_out0[91]),
	.c2v_parallelOut_911(c2v_out1[91]),
	.c2v_parallelOut_912(c2v_out2[91]),
	.c2v_parallelOut_920(c2v_out0[92]),
	.c2v_parallelOut_921(c2v_out1[92]),
	.c2v_parallelOut_922(c2v_out2[92]),
	.c2v_parallelOut_930(c2v_out0[93]),
	.c2v_parallelOut_931(c2v_out1[93]),
	.c2v_parallelOut_932(c2v_out2[93]),
	.c2v_parallelOut_940(c2v_out0[94]),
	.c2v_parallelOut_941(c2v_out1[94]),
	.c2v_parallelOut_942(c2v_out2[94]),
	.c2v_parallelOut_950(c2v_out0[95]),
	.c2v_parallelOut_951(c2v_out1[95]),
	.c2v_parallelOut_952(c2v_out2[95]),
	.c2v_parallelOut_960(c2v_out0[96]),
	.c2v_parallelOut_961(c2v_out1[96]),
	.c2v_parallelOut_962(c2v_out2[96]),
	.c2v_parallelOut_970(c2v_out0[97]),
	.c2v_parallelOut_971(c2v_out1[97]),
	.c2v_parallelOut_972(c2v_out2[97]),
	.c2v_parallelOut_980(c2v_out0[98]),
	.c2v_parallelOut_981(c2v_out1[98]),
	.c2v_parallelOut_982(c2v_out2[98]),
	.c2v_parallelOut_990(c2v_out0[99]),
	.c2v_parallelOut_991(c2v_out1[99]),
	.c2v_parallelOut_992(c2v_out2[99]),
	.c2v_parallelOut_1000(c2v_out0[100]),
	.c2v_parallelOut_1001(c2v_out1[100]),
	.c2v_parallelOut_1002(c2v_out2[100]),
	.c2v_parallelOut_1010(c2v_out0[101]),
	.c2v_parallelOut_1011(c2v_out1[101]),
	.c2v_parallelOut_1012(c2v_out2[101]),
	.c2v_parallelOut_1020(c2v_out0[102]),
	.c2v_parallelOut_1021(c2v_out1[102]),
	.c2v_parallelOut_1022(c2v_out2[102]),
	.c2v_parallelOut_1030(c2v_out0[103]),
	.c2v_parallelOut_1031(c2v_out1[103]),
	.c2v_parallelOut_1032(c2v_out2[103]),
	.c2v_parallelOut_1040(c2v_out0[104]),
	.c2v_parallelOut_1041(c2v_out1[104]),
	.c2v_parallelOut_1042(c2v_out2[104]),
	.c2v_parallelOut_1050(c2v_out0[105]),
	.c2v_parallelOut_1051(c2v_out1[105]),
	.c2v_parallelOut_1052(c2v_out2[105]),
	.c2v_parallelOut_1060(c2v_out0[106]),
	.c2v_parallelOut_1061(c2v_out1[106]),
	.c2v_parallelOut_1062(c2v_out2[106]),
	.c2v_parallelOut_1070(c2v_out0[107]),
	.c2v_parallelOut_1071(c2v_out1[107]),
	.c2v_parallelOut_1072(c2v_out2[107]),
	.c2v_parallelOut_1080(c2v_out0[108]),
	.c2v_parallelOut_1081(c2v_out1[108]),
	.c2v_parallelOut_1082(c2v_out2[108]),
	.c2v_parallelOut_1090(c2v_out0[109]),
	.c2v_parallelOut_1091(c2v_out1[109]),
	.c2v_parallelOut_1092(c2v_out2[109]),
	.c2v_parallelOut_1100(c2v_out0[110]),
	.c2v_parallelOut_1101(c2v_out1[110]),
	.c2v_parallelOut_1102(c2v_out2[110]),
	.c2v_parallelOut_1110(c2v_out0[111]),
	.c2v_parallelOut_1111(c2v_out1[111]),
	.c2v_parallelOut_1112(c2v_out2[111]),
	.c2v_parallelOut_1120(c2v_out0[112]),
	.c2v_parallelOut_1121(c2v_out1[112]),
	.c2v_parallelOut_1122(c2v_out2[112]),
	.c2v_parallelOut_1130(c2v_out0[113]),
	.c2v_parallelOut_1131(c2v_out1[113]),
	.c2v_parallelOut_1132(c2v_out2[113]),
	.c2v_parallelOut_1140(c2v_out0[114]),
	.c2v_parallelOut_1141(c2v_out1[114]),
	.c2v_parallelOut_1142(c2v_out2[114]),
	.c2v_parallelOut_1150(c2v_out0[115]),
	.c2v_parallelOut_1151(c2v_out1[115]),
	.c2v_parallelOut_1152(c2v_out2[115]),
	.c2v_parallelOut_1160(c2v_out0[116]),
	.c2v_parallelOut_1161(c2v_out1[116]),
	.c2v_parallelOut_1162(c2v_out2[116]),
	.c2v_parallelOut_1170(c2v_out0[117]),
	.c2v_parallelOut_1171(c2v_out1[117]),
	.c2v_parallelOut_1172(c2v_out2[117]),
	.c2v_parallelOut_1180(c2v_out0[118]),
	.c2v_parallelOut_1181(c2v_out1[118]),
	.c2v_parallelOut_1182(c2v_out2[118]),
	.c2v_parallelOut_1190(c2v_out0[119]),
	.c2v_parallelOut_1191(c2v_out1[119]),
	.c2v_parallelOut_1192(c2v_out2[119]),
	.c2v_parallelOut_1200(c2v_out0[120]),
	.c2v_parallelOut_1201(c2v_out1[120]),
	.c2v_parallelOut_1202(c2v_out2[120]),
	.c2v_parallelOut_1210(c2v_out0[121]),
	.c2v_parallelOut_1211(c2v_out1[121]),
	.c2v_parallelOut_1212(c2v_out2[121]),
	.c2v_parallelOut_1220(c2v_out0[122]),
	.c2v_parallelOut_1221(c2v_out1[122]),
	.c2v_parallelOut_1222(c2v_out2[122]),
	.c2v_parallelOut_1230(c2v_out0[123]),
	.c2v_parallelOut_1231(c2v_out1[123]),
	.c2v_parallelOut_1232(c2v_out2[123]),
	.c2v_parallelOut_1240(c2v_out0[124]),
	.c2v_parallelOut_1241(c2v_out1[124]),
	.c2v_parallelOut_1242(c2v_out2[124]),
	.c2v_parallelOut_1250(c2v_out0[125]),
	.c2v_parallelOut_1251(c2v_out1[125]),
	.c2v_parallelOut_1252(c2v_out2[125]),
	.c2v_parallelOut_1260(c2v_out0[126]),
	.c2v_parallelOut_1261(c2v_out1[126]),
	.c2v_parallelOut_1262(c2v_out2[126]),
	.c2v_parallelOut_1270(c2v_out0[127]),
	.c2v_parallelOut_1271(c2v_out1[127]),
	.c2v_parallelOut_1272(c2v_out2[127]),
	.c2v_parallelOut_1280(c2v_out0[128]),
	.c2v_parallelOut_1281(c2v_out1[128]),
	.c2v_parallelOut_1282(c2v_out2[128]),
	.c2v_parallelOut_1290(c2v_out0[129]),
	.c2v_parallelOut_1291(c2v_out1[129]),
	.c2v_parallelOut_1292(c2v_out2[129]),
	.c2v_parallelOut_1300(c2v_out0[130]),
	.c2v_parallelOut_1301(c2v_out1[130]),
	.c2v_parallelOut_1302(c2v_out2[130]),
	.c2v_parallelOut_1310(c2v_out0[131]),
	.c2v_parallelOut_1311(c2v_out1[131]),
	.c2v_parallelOut_1312(c2v_out2[131]),
	.c2v_parallelOut_1320(c2v_out0[132]),
	.c2v_parallelOut_1321(c2v_out1[132]),
	.c2v_parallelOut_1322(c2v_out2[132]),
	.c2v_parallelOut_1330(c2v_out0[133]),
	.c2v_parallelOut_1331(c2v_out1[133]),
	.c2v_parallelOut_1332(c2v_out2[133]),
	.c2v_parallelOut_1340(c2v_out0[134]),
	.c2v_parallelOut_1341(c2v_out1[134]),
	.c2v_parallelOut_1342(c2v_out2[134]),
	.c2v_parallelOut_1350(c2v_out0[135]),
	.c2v_parallelOut_1351(c2v_out1[135]),
	.c2v_parallelOut_1352(c2v_out2[135]),
	.c2v_parallelOut_1360(c2v_out0[136]),
	.c2v_parallelOut_1361(c2v_out1[136]),
	.c2v_parallelOut_1362(c2v_out2[136]),
	.c2v_parallelOut_1370(c2v_out0[137]),
	.c2v_parallelOut_1371(c2v_out1[137]),
	.c2v_parallelOut_1372(c2v_out2[137]),
	.c2v_parallelOut_1380(c2v_out0[138]),
	.c2v_parallelOut_1381(c2v_out1[138]),
	.c2v_parallelOut_1382(c2v_out2[138]),
	.c2v_parallelOut_1390(c2v_out0[139]),
	.c2v_parallelOut_1391(c2v_out1[139]),
	.c2v_parallelOut_1392(c2v_out2[139]),
	.c2v_parallelOut_1400(c2v_out0[140]),
	.c2v_parallelOut_1401(c2v_out1[140]),
	.c2v_parallelOut_1402(c2v_out2[140]),
	.c2v_parallelOut_1410(c2v_out0[141]),
	.c2v_parallelOut_1411(c2v_out1[141]),
	.c2v_parallelOut_1412(c2v_out2[141]),
	.c2v_parallelOut_1420(c2v_out0[142]),
	.c2v_parallelOut_1421(c2v_out1[142]),
	.c2v_parallelOut_1422(c2v_out2[142]),
	.c2v_parallelOut_1430(c2v_out0[143]),
	.c2v_parallelOut_1431(c2v_out1[143]),
	.c2v_parallelOut_1432(c2v_out2[143]),
	.c2v_parallelOut_1440(c2v_out0[144]),
	.c2v_parallelOut_1441(c2v_out1[144]),
	.c2v_parallelOut_1442(c2v_out2[144]),
	.c2v_parallelOut_1450(c2v_out0[145]),
	.c2v_parallelOut_1451(c2v_out1[145]),
	.c2v_parallelOut_1452(c2v_out2[145]),
	.c2v_parallelOut_1460(c2v_out0[146]),
	.c2v_parallelOut_1461(c2v_out1[146]),
	.c2v_parallelOut_1462(c2v_out2[146]),
	.c2v_parallelOut_1470(c2v_out0[147]),
	.c2v_parallelOut_1471(c2v_out1[147]),
	.c2v_parallelOut_1472(c2v_out2[147]),
	.c2v_parallelOut_1480(c2v_out0[148]),
	.c2v_parallelOut_1481(c2v_out1[148]),
	.c2v_parallelOut_1482(c2v_out2[148]),
	.c2v_parallelOut_1490(c2v_out0[149]),
	.c2v_parallelOut_1491(c2v_out1[149]),
	.c2v_parallelOut_1492(c2v_out2[149]),
	.c2v_parallelOut_1500(c2v_out0[150]),
	.c2v_parallelOut_1501(c2v_out1[150]),
	.c2v_parallelOut_1502(c2v_out2[150]),
	.c2v_parallelOut_1510(c2v_out0[151]),
	.c2v_parallelOut_1511(c2v_out1[151]),
	.c2v_parallelOut_1512(c2v_out2[151]),
	.c2v_parallelOut_1520(c2v_out0[152]),
	.c2v_parallelOut_1521(c2v_out1[152]),
	.c2v_parallelOut_1522(c2v_out2[152]),
	.c2v_parallelOut_1530(c2v_out0[153]),
	.c2v_parallelOut_1531(c2v_out1[153]),
	.c2v_parallelOut_1532(c2v_out2[153]),
	.c2v_parallelOut_1540(c2v_out0[154]),
	.c2v_parallelOut_1541(c2v_out1[154]),
	.c2v_parallelOut_1542(c2v_out2[154]),
	.c2v_parallelOut_1550(c2v_out0[155]),
	.c2v_parallelOut_1551(c2v_out1[155]),
	.c2v_parallelOut_1552(c2v_out2[155]),
	.c2v_parallelOut_1560(c2v_out0[156]),
	.c2v_parallelOut_1561(c2v_out1[156]),
	.c2v_parallelOut_1562(c2v_out2[156]),
	.c2v_parallelOut_1570(c2v_out0[157]),
	.c2v_parallelOut_1571(c2v_out1[157]),
	.c2v_parallelOut_1572(c2v_out2[157]),
	.c2v_parallelOut_1580(c2v_out0[158]),
	.c2v_parallelOut_1581(c2v_out1[158]),
	.c2v_parallelOut_1582(c2v_out2[158]),
	.c2v_parallelOut_1590(c2v_out0[159]),
	.c2v_parallelOut_1591(c2v_out1[159]),
	.c2v_parallelOut_1592(c2v_out2[159]),
	.c2v_parallelOut_1600(c2v_out0[160]),
	.c2v_parallelOut_1601(c2v_out1[160]),
	.c2v_parallelOut_1602(c2v_out2[160]),
	.c2v_parallelOut_1610(c2v_out0[161]),
	.c2v_parallelOut_1611(c2v_out1[161]),
	.c2v_parallelOut_1612(c2v_out2[161]),
	.c2v_parallelOut_1620(c2v_out0[162]),
	.c2v_parallelOut_1621(c2v_out1[162]),
	.c2v_parallelOut_1622(c2v_out2[162]),
	.c2v_parallelOut_1630(c2v_out0[163]),
	.c2v_parallelOut_1631(c2v_out1[163]),
	.c2v_parallelOut_1632(c2v_out2[163]),
	.c2v_parallelOut_1640(c2v_out0[164]),
	.c2v_parallelOut_1641(c2v_out1[164]),
	.c2v_parallelOut_1642(c2v_out2[164]),
	.c2v_parallelOut_1650(c2v_out0[165]),
	.c2v_parallelOut_1651(c2v_out1[165]),
	.c2v_parallelOut_1652(c2v_out2[165]),
	.c2v_parallelOut_1660(c2v_out0[166]),
	.c2v_parallelOut_1661(c2v_out1[166]),
	.c2v_parallelOut_1662(c2v_out2[166]),
	.c2v_parallelOut_1670(c2v_out0[167]),
	.c2v_parallelOut_1671(c2v_out1[167]),
	.c2v_parallelOut_1672(c2v_out2[167]),
	.c2v_parallelOut_1680(c2v_out0[168]),
	.c2v_parallelOut_1681(c2v_out1[168]),
	.c2v_parallelOut_1682(c2v_out2[168]),
	.c2v_parallelOut_1690(c2v_out0[169]),
	.c2v_parallelOut_1691(c2v_out1[169]),
	.c2v_parallelOut_1692(c2v_out2[169]),
	.c2v_parallelOut_1700(c2v_out0[170]),
	.c2v_parallelOut_1701(c2v_out1[170]),
	.c2v_parallelOut_1702(c2v_out2[170]),
	.c2v_parallelOut_1710(c2v_out0[171]),
	.c2v_parallelOut_1711(c2v_out1[171]),
	.c2v_parallelOut_1712(c2v_out2[171]),
	.c2v_parallelOut_1720(c2v_out0[172]),
	.c2v_parallelOut_1721(c2v_out1[172]),
	.c2v_parallelOut_1722(c2v_out2[172]),
	.c2v_parallelOut_1730(c2v_out0[173]),
	.c2v_parallelOut_1731(c2v_out1[173]),
	.c2v_parallelOut_1732(c2v_out2[173]),
	.c2v_parallelOut_1740(c2v_out0[174]),
	.c2v_parallelOut_1741(c2v_out1[174]),
	.c2v_parallelOut_1742(c2v_out2[174]),
	.c2v_parallelOut_1750(c2v_out0[175]),
	.c2v_parallelOut_1751(c2v_out1[175]),
	.c2v_parallelOut_1752(c2v_out2[175]),
	.c2v_parallelOut_1760(c2v_out0[176]),
	.c2v_parallelOut_1761(c2v_out1[176]),
	.c2v_parallelOut_1762(c2v_out2[176]),
	.c2v_parallelOut_1770(c2v_out0[177]),
	.c2v_parallelOut_1771(c2v_out1[177]),
	.c2v_parallelOut_1772(c2v_out2[177]),
	.c2v_parallelOut_1780(c2v_out0[178]),
	.c2v_parallelOut_1781(c2v_out1[178]),
	.c2v_parallelOut_1782(c2v_out2[178]),
	.c2v_parallelOut_1790(c2v_out0[179]),
	.c2v_parallelOut_1791(c2v_out1[179]),
	.c2v_parallelOut_1792(c2v_out2[179]),
	.c2v_parallelOut_1800(c2v_out0[180]),
	.c2v_parallelOut_1801(c2v_out1[180]),
	.c2v_parallelOut_1802(c2v_out2[180]),
	.c2v_parallelOut_1810(c2v_out0[181]),
	.c2v_parallelOut_1811(c2v_out1[181]),
	.c2v_parallelOut_1812(c2v_out2[181]),
	.c2v_parallelOut_1820(c2v_out0[182]),
	.c2v_parallelOut_1821(c2v_out1[182]),
	.c2v_parallelOut_1822(c2v_out2[182]),
	.c2v_parallelOut_1830(c2v_out0[183]),
	.c2v_parallelOut_1831(c2v_out1[183]),
	.c2v_parallelOut_1832(c2v_out2[183]),
	.c2v_parallelOut_1840(c2v_out0[184]),
	.c2v_parallelOut_1841(c2v_out1[184]),
	.c2v_parallelOut_1842(c2v_out2[184]),
	.c2v_parallelOut_1850(c2v_out0[185]),
	.c2v_parallelOut_1851(c2v_out1[185]),
	.c2v_parallelOut_1852(c2v_out2[185]),
	.c2v_parallelOut_1860(c2v_out0[186]),
	.c2v_parallelOut_1861(c2v_out1[186]),
	.c2v_parallelOut_1862(c2v_out2[186]),
	.c2v_parallelOut_1870(c2v_out0[187]),
	.c2v_parallelOut_1871(c2v_out1[187]),
	.c2v_parallelOut_1872(c2v_out2[187]),
	.c2v_parallelOut_1880(c2v_out0[188]),
	.c2v_parallelOut_1881(c2v_out1[188]),
	.c2v_parallelOut_1882(c2v_out2[188]),
	.c2v_parallelOut_1890(c2v_out0[189]),
	.c2v_parallelOut_1891(c2v_out1[189]),
	.c2v_parallelOut_1892(c2v_out2[189]),
	.c2v_parallelOut_1900(c2v_out0[190]),
	.c2v_parallelOut_1901(c2v_out1[190]),
	.c2v_parallelOut_1902(c2v_out2[190]),
	.c2v_parallelOut_1910(c2v_out0[191]),
	.c2v_parallelOut_1911(c2v_out1[191]),
	.c2v_parallelOut_1912(c2v_out2[191]),
	.c2v_parallelOut_1920(c2v_out0[192]),
	.c2v_parallelOut_1921(c2v_out1[192]),
	.c2v_parallelOut_1922(c2v_out2[192]),
	.c2v_parallelOut_1930(c2v_out0[193]),
	.c2v_parallelOut_1931(c2v_out1[193]),
	.c2v_parallelOut_1932(c2v_out2[193]),
	.c2v_parallelOut_1940(c2v_out0[194]),
	.c2v_parallelOut_1941(c2v_out1[194]),
	.c2v_parallelOut_1942(c2v_out2[194]),
	.c2v_parallelOut_1950(c2v_out0[195]),
	.c2v_parallelOut_1951(c2v_out1[195]),
	.c2v_parallelOut_1952(c2v_out2[195]),
	.c2v_parallelOut_1960(c2v_out0[196]),
	.c2v_parallelOut_1961(c2v_out1[196]),
	.c2v_parallelOut_1962(c2v_out2[196]),
	.c2v_parallelOut_1970(c2v_out0[197]),
	.c2v_parallelOut_1971(c2v_out1[197]),
	.c2v_parallelOut_1972(c2v_out2[197]),
	.c2v_parallelOut_1980(c2v_out0[198]),
	.c2v_parallelOut_1981(c2v_out1[198]),
	.c2v_parallelOut_1982(c2v_out2[198]),
	.c2v_parallelOut_1990(c2v_out0[199]),
	.c2v_parallelOut_1991(c2v_out1[199]),
	.c2v_parallelOut_1992(c2v_out2[199]),
	.c2v_parallelOut_2000(c2v_out0[200]),
	.c2v_parallelOut_2001(c2v_out1[200]),
	.c2v_parallelOut_2002(c2v_out2[200]),
	.c2v_parallelOut_2010(c2v_out0[201]),
	.c2v_parallelOut_2011(c2v_out1[201]),
	.c2v_parallelOut_2012(c2v_out2[201]),
	.c2v_parallelOut_2020(c2v_out0[202]),
	.c2v_parallelOut_2021(c2v_out1[202]),
	.c2v_parallelOut_2022(c2v_out2[202]),
	.c2v_parallelOut_2030(c2v_out0[203]),
	.c2v_parallelOut_2031(c2v_out1[203]),
	.c2v_parallelOut_2032(c2v_out2[203]),
	
	.c2v_parallelIn_00(c2v_0[0]),
	.c2v_parallelIn_01(c2v_1[0]),
	.c2v_parallelIn_02(c2v_2[0]),
	.c2v_parallelIn_03(c2v_3[0]),
	.c2v_parallelIn_04(c2v_4[0]),
	.c2v_parallelIn_05(c2v_5[0]),
	.c2v_parallelIn_10(c2v_0[1]),
	.c2v_parallelIn_11(c2v_1[1]),
	.c2v_parallelIn_12(c2v_2[1]),
	.c2v_parallelIn_13(c2v_3[1]),
	.c2v_parallelIn_14(c2v_4[1]),
	.c2v_parallelIn_15(c2v_5[1]),
	.c2v_parallelIn_20(c2v_0[2]),
	.c2v_parallelIn_21(c2v_1[2]),
	.c2v_parallelIn_22(c2v_2[2]),
	.c2v_parallelIn_23(c2v_3[2]),
	.c2v_parallelIn_24(c2v_4[2]),
	.c2v_parallelIn_25(c2v_5[2]),
	.c2v_parallelIn_30(c2v_0[3]),
	.c2v_parallelIn_31(c2v_1[3]),
	.c2v_parallelIn_32(c2v_2[3]),
	.c2v_parallelIn_33(c2v_3[3]),
	.c2v_parallelIn_34(c2v_4[3]),
	.c2v_parallelIn_35(c2v_5[3]),
	.c2v_parallelIn_40(c2v_0[4]),
	.c2v_parallelIn_41(c2v_1[4]),
	.c2v_parallelIn_42(c2v_2[4]),
	.c2v_parallelIn_43(c2v_3[4]),
	.c2v_parallelIn_44(c2v_4[4]),
	.c2v_parallelIn_45(c2v_5[4]),
	.c2v_parallelIn_50(c2v_0[5]),
	.c2v_parallelIn_51(c2v_1[5]),
	.c2v_parallelIn_52(c2v_2[5]),
	.c2v_parallelIn_53(c2v_3[5]),
	.c2v_parallelIn_54(c2v_4[5]),
	.c2v_parallelIn_55(c2v_5[5]),
	.c2v_parallelIn_60(c2v_0[6]),
	.c2v_parallelIn_61(c2v_1[6]),
	.c2v_parallelIn_62(c2v_2[6]),
	.c2v_parallelIn_63(c2v_3[6]),
	.c2v_parallelIn_64(c2v_4[6]),
	.c2v_parallelIn_65(c2v_5[6]),
	.c2v_parallelIn_70(c2v_0[7]),
	.c2v_parallelIn_71(c2v_1[7]),
	.c2v_parallelIn_72(c2v_2[7]),
	.c2v_parallelIn_73(c2v_3[7]),
	.c2v_parallelIn_74(c2v_4[7]),
	.c2v_parallelIn_75(c2v_5[7]),
	.c2v_parallelIn_80(c2v_0[8]),
	.c2v_parallelIn_81(c2v_1[8]),
	.c2v_parallelIn_82(c2v_2[8]),
	.c2v_parallelIn_83(c2v_3[8]),
	.c2v_parallelIn_84(c2v_4[8]),
	.c2v_parallelIn_85(c2v_5[8]),
	.c2v_parallelIn_90(c2v_0[9]),
	.c2v_parallelIn_91(c2v_1[9]),
	.c2v_parallelIn_92(c2v_2[9]),
	.c2v_parallelIn_93(c2v_3[9]),
	.c2v_parallelIn_94(c2v_4[9]),
	.c2v_parallelIn_95(c2v_5[9]),
	.c2v_parallelIn_100(c2v_0[10]),
	.c2v_parallelIn_101(c2v_1[10]),
	.c2v_parallelIn_102(c2v_2[10]),
	.c2v_parallelIn_103(c2v_3[10]),
	.c2v_parallelIn_104(c2v_4[10]),
	.c2v_parallelIn_105(c2v_5[10]),
	.c2v_parallelIn_110(c2v_0[11]),
	.c2v_parallelIn_111(c2v_1[11]),
	.c2v_parallelIn_112(c2v_2[11]),
	.c2v_parallelIn_113(c2v_3[11]),
	.c2v_parallelIn_114(c2v_4[11]),
	.c2v_parallelIn_115(c2v_5[11]),
	.c2v_parallelIn_120(c2v_0[12]),
	.c2v_parallelIn_121(c2v_1[12]),
	.c2v_parallelIn_122(c2v_2[12]),
	.c2v_parallelIn_123(c2v_3[12]),
	.c2v_parallelIn_124(c2v_4[12]),
	.c2v_parallelIn_125(c2v_5[12]),
	.c2v_parallelIn_130(c2v_0[13]),
	.c2v_parallelIn_131(c2v_1[13]),
	.c2v_parallelIn_132(c2v_2[13]),
	.c2v_parallelIn_133(c2v_3[13]),
	.c2v_parallelIn_134(c2v_4[13]),
	.c2v_parallelIn_135(c2v_5[13]),
	.c2v_parallelIn_140(c2v_0[14]),
	.c2v_parallelIn_141(c2v_1[14]),
	.c2v_parallelIn_142(c2v_2[14]),
	.c2v_parallelIn_143(c2v_3[14]),
	.c2v_parallelIn_144(c2v_4[14]),
	.c2v_parallelIn_145(c2v_5[14]),
	.c2v_parallelIn_150(c2v_0[15]),
	.c2v_parallelIn_151(c2v_1[15]),
	.c2v_parallelIn_152(c2v_2[15]),
	.c2v_parallelIn_153(c2v_3[15]),
	.c2v_parallelIn_154(c2v_4[15]),
	.c2v_parallelIn_155(c2v_5[15]),
	.c2v_parallelIn_160(c2v_0[16]),
	.c2v_parallelIn_161(c2v_1[16]),
	.c2v_parallelIn_162(c2v_2[16]),
	.c2v_parallelIn_163(c2v_3[16]),
	.c2v_parallelIn_164(c2v_4[16]),
	.c2v_parallelIn_165(c2v_5[16]),
	.c2v_parallelIn_170(c2v_0[17]),
	.c2v_parallelIn_171(c2v_1[17]),
	.c2v_parallelIn_172(c2v_2[17]),
	.c2v_parallelIn_173(c2v_3[17]),
	.c2v_parallelIn_174(c2v_4[17]),
	.c2v_parallelIn_175(c2v_5[17]),
	.c2v_parallelIn_180(c2v_0[18]),
	.c2v_parallelIn_181(c2v_1[18]),
	.c2v_parallelIn_182(c2v_2[18]),
	.c2v_parallelIn_183(c2v_3[18]),
	.c2v_parallelIn_184(c2v_4[18]),
	.c2v_parallelIn_185(c2v_5[18]),
	.c2v_parallelIn_190(c2v_0[19]),
	.c2v_parallelIn_191(c2v_1[19]),
	.c2v_parallelIn_192(c2v_2[19]),
	.c2v_parallelIn_193(c2v_3[19]),
	.c2v_parallelIn_194(c2v_4[19]),
	.c2v_parallelIn_195(c2v_5[19]),
	.c2v_parallelIn_200(c2v_0[20]),
	.c2v_parallelIn_201(c2v_1[20]),
	.c2v_parallelIn_202(c2v_2[20]),
	.c2v_parallelIn_203(c2v_3[20]),
	.c2v_parallelIn_204(c2v_4[20]),
	.c2v_parallelIn_205(c2v_5[20]),
	.c2v_parallelIn_210(c2v_0[21]),
	.c2v_parallelIn_211(c2v_1[21]),
	.c2v_parallelIn_212(c2v_2[21]),
	.c2v_parallelIn_213(c2v_3[21]),
	.c2v_parallelIn_214(c2v_4[21]),
	.c2v_parallelIn_215(c2v_5[21]),
	.c2v_parallelIn_220(c2v_0[22]),
	.c2v_parallelIn_221(c2v_1[22]),
	.c2v_parallelIn_222(c2v_2[22]),
	.c2v_parallelIn_223(c2v_3[22]),
	.c2v_parallelIn_224(c2v_4[22]),
	.c2v_parallelIn_225(c2v_5[22]),
	.c2v_parallelIn_230(c2v_0[23]),
	.c2v_parallelIn_231(c2v_1[23]),
	.c2v_parallelIn_232(c2v_2[23]),
	.c2v_parallelIn_233(c2v_3[23]),
	.c2v_parallelIn_234(c2v_4[23]),
	.c2v_parallelIn_235(c2v_5[23]),
	.c2v_parallelIn_240(c2v_0[24]),
	.c2v_parallelIn_241(c2v_1[24]),
	.c2v_parallelIn_242(c2v_2[24]),
	.c2v_parallelIn_243(c2v_3[24]),
	.c2v_parallelIn_244(c2v_4[24]),
	.c2v_parallelIn_245(c2v_5[24]),
	.c2v_parallelIn_250(c2v_0[25]),
	.c2v_parallelIn_251(c2v_1[25]),
	.c2v_parallelIn_252(c2v_2[25]),
	.c2v_parallelIn_253(c2v_3[25]),
	.c2v_parallelIn_254(c2v_4[25]),
	.c2v_parallelIn_255(c2v_5[25]),
	.c2v_parallelIn_260(c2v_0[26]),
	.c2v_parallelIn_261(c2v_1[26]),
	.c2v_parallelIn_262(c2v_2[26]),
	.c2v_parallelIn_263(c2v_3[26]),
	.c2v_parallelIn_264(c2v_4[26]),
	.c2v_parallelIn_265(c2v_5[26]),
	.c2v_parallelIn_270(c2v_0[27]),
	.c2v_parallelIn_271(c2v_1[27]),
	.c2v_parallelIn_272(c2v_2[27]),
	.c2v_parallelIn_273(c2v_3[27]),
	.c2v_parallelIn_274(c2v_4[27]),
	.c2v_parallelIn_275(c2v_5[27]),
	.c2v_parallelIn_280(c2v_0[28]),
	.c2v_parallelIn_281(c2v_1[28]),
	.c2v_parallelIn_282(c2v_2[28]),
	.c2v_parallelIn_283(c2v_3[28]),
	.c2v_parallelIn_284(c2v_4[28]),
	.c2v_parallelIn_285(c2v_5[28]),
	.c2v_parallelIn_290(c2v_0[29]),
	.c2v_parallelIn_291(c2v_1[29]),
	.c2v_parallelIn_292(c2v_2[29]),
	.c2v_parallelIn_293(c2v_3[29]),
	.c2v_parallelIn_294(c2v_4[29]),
	.c2v_parallelIn_295(c2v_5[29]),
	.c2v_parallelIn_300(c2v_0[30]),
	.c2v_parallelIn_301(c2v_1[30]),
	.c2v_parallelIn_302(c2v_2[30]),
	.c2v_parallelIn_303(c2v_3[30]),
	.c2v_parallelIn_304(c2v_4[30]),
	.c2v_parallelIn_305(c2v_5[30]),
	.c2v_parallelIn_310(c2v_0[31]),
	.c2v_parallelIn_311(c2v_1[31]),
	.c2v_parallelIn_312(c2v_2[31]),
	.c2v_parallelIn_313(c2v_3[31]),
	.c2v_parallelIn_314(c2v_4[31]),
	.c2v_parallelIn_315(c2v_5[31]),
	.c2v_parallelIn_320(c2v_0[32]),
	.c2v_parallelIn_321(c2v_1[32]),
	.c2v_parallelIn_322(c2v_2[32]),
	.c2v_parallelIn_323(c2v_3[32]),
	.c2v_parallelIn_324(c2v_4[32]),
	.c2v_parallelIn_325(c2v_5[32]),
	.c2v_parallelIn_330(c2v_0[33]),
	.c2v_parallelIn_331(c2v_1[33]),
	.c2v_parallelIn_332(c2v_2[33]),
	.c2v_parallelIn_333(c2v_3[33]),
	.c2v_parallelIn_334(c2v_4[33]),
	.c2v_parallelIn_335(c2v_5[33]),
	.c2v_parallelIn_340(c2v_0[34]),
	.c2v_parallelIn_341(c2v_1[34]),
	.c2v_parallelIn_342(c2v_2[34]),
	.c2v_parallelIn_343(c2v_3[34]),
	.c2v_parallelIn_344(c2v_4[34]),
	.c2v_parallelIn_345(c2v_5[34]),
	.c2v_parallelIn_350(c2v_0[35]),
	.c2v_parallelIn_351(c2v_1[35]),
	.c2v_parallelIn_352(c2v_2[35]),
	.c2v_parallelIn_353(c2v_3[35]),
	.c2v_parallelIn_354(c2v_4[35]),
	.c2v_parallelIn_355(c2v_5[35]),
	.c2v_parallelIn_360(c2v_0[36]),
	.c2v_parallelIn_361(c2v_1[36]),
	.c2v_parallelIn_362(c2v_2[36]),
	.c2v_parallelIn_363(c2v_3[36]),
	.c2v_parallelIn_364(c2v_4[36]),
	.c2v_parallelIn_365(c2v_5[36]),
	.c2v_parallelIn_370(c2v_0[37]),
	.c2v_parallelIn_371(c2v_1[37]),
	.c2v_parallelIn_372(c2v_2[37]),
	.c2v_parallelIn_373(c2v_3[37]),
	.c2v_parallelIn_374(c2v_4[37]),
	.c2v_parallelIn_375(c2v_5[37]),
	.c2v_parallelIn_380(c2v_0[38]),
	.c2v_parallelIn_381(c2v_1[38]),
	.c2v_parallelIn_382(c2v_2[38]),
	.c2v_parallelIn_383(c2v_3[38]),
	.c2v_parallelIn_384(c2v_4[38]),
	.c2v_parallelIn_385(c2v_5[38]),
	.c2v_parallelIn_390(c2v_0[39]),
	.c2v_parallelIn_391(c2v_1[39]),
	.c2v_parallelIn_392(c2v_2[39]),
	.c2v_parallelIn_393(c2v_3[39]),
	.c2v_parallelIn_394(c2v_4[39]),
	.c2v_parallelIn_395(c2v_5[39]),
	.c2v_parallelIn_400(c2v_0[40]),
	.c2v_parallelIn_401(c2v_1[40]),
	.c2v_parallelIn_402(c2v_2[40]),
	.c2v_parallelIn_403(c2v_3[40]),
	.c2v_parallelIn_404(c2v_4[40]),
	.c2v_parallelIn_405(c2v_5[40]),
	.c2v_parallelIn_410(c2v_0[41]),
	.c2v_parallelIn_411(c2v_1[41]),
	.c2v_parallelIn_412(c2v_2[41]),
	.c2v_parallelIn_413(c2v_3[41]),
	.c2v_parallelIn_414(c2v_4[41]),
	.c2v_parallelIn_415(c2v_5[41]),
	.c2v_parallelIn_420(c2v_0[42]),
	.c2v_parallelIn_421(c2v_1[42]),
	.c2v_parallelIn_422(c2v_2[42]),
	.c2v_parallelIn_423(c2v_3[42]),
	.c2v_parallelIn_424(c2v_4[42]),
	.c2v_parallelIn_425(c2v_5[42]),
	.c2v_parallelIn_430(c2v_0[43]),
	.c2v_parallelIn_431(c2v_1[43]),
	.c2v_parallelIn_432(c2v_2[43]),
	.c2v_parallelIn_433(c2v_3[43]),
	.c2v_parallelIn_434(c2v_4[43]),
	.c2v_parallelIn_435(c2v_5[43]),
	.c2v_parallelIn_440(c2v_0[44]),
	.c2v_parallelIn_441(c2v_1[44]),
	.c2v_parallelIn_442(c2v_2[44]),
	.c2v_parallelIn_443(c2v_3[44]),
	.c2v_parallelIn_444(c2v_4[44]),
	.c2v_parallelIn_445(c2v_5[44]),
	.c2v_parallelIn_450(c2v_0[45]),
	.c2v_parallelIn_451(c2v_1[45]),
	.c2v_parallelIn_452(c2v_2[45]),
	.c2v_parallelIn_453(c2v_3[45]),
	.c2v_parallelIn_454(c2v_4[45]),
	.c2v_parallelIn_455(c2v_5[45]),
	.c2v_parallelIn_460(c2v_0[46]),
	.c2v_parallelIn_461(c2v_1[46]),
	.c2v_parallelIn_462(c2v_2[46]),
	.c2v_parallelIn_463(c2v_3[46]),
	.c2v_parallelIn_464(c2v_4[46]),
	.c2v_parallelIn_465(c2v_5[46]),
	.c2v_parallelIn_470(c2v_0[47]),
	.c2v_parallelIn_471(c2v_1[47]),
	.c2v_parallelIn_472(c2v_2[47]),
	.c2v_parallelIn_473(c2v_3[47]),
	.c2v_parallelIn_474(c2v_4[47]),
	.c2v_parallelIn_475(c2v_5[47]),
	.c2v_parallelIn_480(c2v_0[48]),
	.c2v_parallelIn_481(c2v_1[48]),
	.c2v_parallelIn_482(c2v_2[48]),
	.c2v_parallelIn_483(c2v_3[48]),
	.c2v_parallelIn_484(c2v_4[48]),
	.c2v_parallelIn_485(c2v_5[48]),
	.c2v_parallelIn_490(c2v_0[49]),
	.c2v_parallelIn_491(c2v_1[49]),
	.c2v_parallelIn_492(c2v_2[49]),
	.c2v_parallelIn_493(c2v_3[49]),
	.c2v_parallelIn_494(c2v_4[49]),
	.c2v_parallelIn_495(c2v_5[49]),
	.c2v_parallelIn_500(c2v_0[50]),
	.c2v_parallelIn_501(c2v_1[50]),
	.c2v_parallelIn_502(c2v_2[50]),
	.c2v_parallelIn_503(c2v_3[50]),
	.c2v_parallelIn_504(c2v_4[50]),
	.c2v_parallelIn_505(c2v_5[50]),
	.c2v_parallelIn_510(c2v_0[51]),
	.c2v_parallelIn_511(c2v_1[51]),
	.c2v_parallelIn_512(c2v_2[51]),
	.c2v_parallelIn_513(c2v_3[51]),
	.c2v_parallelIn_514(c2v_4[51]),
	.c2v_parallelIn_515(c2v_5[51]),
	.c2v_parallelIn_520(c2v_0[52]),
	.c2v_parallelIn_521(c2v_1[52]),
	.c2v_parallelIn_522(c2v_2[52]),
	.c2v_parallelIn_523(c2v_3[52]),
	.c2v_parallelIn_524(c2v_4[52]),
	.c2v_parallelIn_525(c2v_5[52]),
	.c2v_parallelIn_530(c2v_0[53]),
	.c2v_parallelIn_531(c2v_1[53]),
	.c2v_parallelIn_532(c2v_2[53]),
	.c2v_parallelIn_533(c2v_3[53]),
	.c2v_parallelIn_534(c2v_4[53]),
	.c2v_parallelIn_535(c2v_5[53]),
	.c2v_parallelIn_540(c2v_0[54]),
	.c2v_parallelIn_541(c2v_1[54]),
	.c2v_parallelIn_542(c2v_2[54]),
	.c2v_parallelIn_543(c2v_3[54]),
	.c2v_parallelIn_544(c2v_4[54]),
	.c2v_parallelIn_545(c2v_5[54]),
	.c2v_parallelIn_550(c2v_0[55]),
	.c2v_parallelIn_551(c2v_1[55]),
	.c2v_parallelIn_552(c2v_2[55]),
	.c2v_parallelIn_553(c2v_3[55]),
	.c2v_parallelIn_554(c2v_4[55]),
	.c2v_parallelIn_555(c2v_5[55]),
	.c2v_parallelIn_560(c2v_0[56]),
	.c2v_parallelIn_561(c2v_1[56]),
	.c2v_parallelIn_562(c2v_2[56]),
	.c2v_parallelIn_563(c2v_3[56]),
	.c2v_parallelIn_564(c2v_4[56]),
	.c2v_parallelIn_565(c2v_5[56]),
	.c2v_parallelIn_570(c2v_0[57]),
	.c2v_parallelIn_571(c2v_1[57]),
	.c2v_parallelIn_572(c2v_2[57]),
	.c2v_parallelIn_573(c2v_3[57]),
	.c2v_parallelIn_574(c2v_4[57]),
	.c2v_parallelIn_575(c2v_5[57]),
	.c2v_parallelIn_580(c2v_0[58]),
	.c2v_parallelIn_581(c2v_1[58]),
	.c2v_parallelIn_582(c2v_2[58]),
	.c2v_parallelIn_583(c2v_3[58]),
	.c2v_parallelIn_584(c2v_4[58]),
	.c2v_parallelIn_585(c2v_5[58]),
	.c2v_parallelIn_590(c2v_0[59]),
	.c2v_parallelIn_591(c2v_1[59]),
	.c2v_parallelIn_592(c2v_2[59]),
	.c2v_parallelIn_593(c2v_3[59]),
	.c2v_parallelIn_594(c2v_4[59]),
	.c2v_parallelIn_595(c2v_5[59]),
	.c2v_parallelIn_600(c2v_0[60]),
	.c2v_parallelIn_601(c2v_1[60]),
	.c2v_parallelIn_602(c2v_2[60]),
	.c2v_parallelIn_603(c2v_3[60]),
	.c2v_parallelIn_604(c2v_4[60]),
	.c2v_parallelIn_605(c2v_5[60]),
	.c2v_parallelIn_610(c2v_0[61]),
	.c2v_parallelIn_611(c2v_1[61]),
	.c2v_parallelIn_612(c2v_2[61]),
	.c2v_parallelIn_613(c2v_3[61]),
	.c2v_parallelIn_614(c2v_4[61]),
	.c2v_parallelIn_615(c2v_5[61]),
	.c2v_parallelIn_620(c2v_0[62]),
	.c2v_parallelIn_621(c2v_1[62]),
	.c2v_parallelIn_622(c2v_2[62]),
	.c2v_parallelIn_623(c2v_3[62]),
	.c2v_parallelIn_624(c2v_4[62]),
	.c2v_parallelIn_625(c2v_5[62]),
	.c2v_parallelIn_630(c2v_0[63]),
	.c2v_parallelIn_631(c2v_1[63]),
	.c2v_parallelIn_632(c2v_2[63]),
	.c2v_parallelIn_633(c2v_3[63]),
	.c2v_parallelIn_634(c2v_4[63]),
	.c2v_parallelIn_635(c2v_5[63]),
	.c2v_parallelIn_640(c2v_0[64]),
	.c2v_parallelIn_641(c2v_1[64]),
	.c2v_parallelIn_642(c2v_2[64]),
	.c2v_parallelIn_643(c2v_3[64]),
	.c2v_parallelIn_644(c2v_4[64]),
	.c2v_parallelIn_645(c2v_5[64]),
	.c2v_parallelIn_650(c2v_0[65]),
	.c2v_parallelIn_651(c2v_1[65]),
	.c2v_parallelIn_652(c2v_2[65]),
	.c2v_parallelIn_653(c2v_3[65]),
	.c2v_parallelIn_654(c2v_4[65]),
	.c2v_parallelIn_655(c2v_5[65]),
	.c2v_parallelIn_660(c2v_0[66]),
	.c2v_parallelIn_661(c2v_1[66]),
	.c2v_parallelIn_662(c2v_2[66]),
	.c2v_parallelIn_663(c2v_3[66]),
	.c2v_parallelIn_664(c2v_4[66]),
	.c2v_parallelIn_665(c2v_5[66]),
	.c2v_parallelIn_670(c2v_0[67]),
	.c2v_parallelIn_671(c2v_1[67]),
	.c2v_parallelIn_672(c2v_2[67]),
	.c2v_parallelIn_673(c2v_3[67]),
	.c2v_parallelIn_674(c2v_4[67]),
	.c2v_parallelIn_675(c2v_5[67]),
	.c2v_parallelIn_680(c2v_0[68]),
	.c2v_parallelIn_681(c2v_1[68]),
	.c2v_parallelIn_682(c2v_2[68]),
	.c2v_parallelIn_683(c2v_3[68]),
	.c2v_parallelIn_684(c2v_4[68]),
	.c2v_parallelIn_685(c2v_5[68]),
	.c2v_parallelIn_690(c2v_0[69]),
	.c2v_parallelIn_691(c2v_1[69]),
	.c2v_parallelIn_692(c2v_2[69]),
	.c2v_parallelIn_693(c2v_3[69]),
	.c2v_parallelIn_694(c2v_4[69]),
	.c2v_parallelIn_695(c2v_5[69]),
	.c2v_parallelIn_700(c2v_0[70]),
	.c2v_parallelIn_701(c2v_1[70]),
	.c2v_parallelIn_702(c2v_2[70]),
	.c2v_parallelIn_703(c2v_3[70]),
	.c2v_parallelIn_704(c2v_4[70]),
	.c2v_parallelIn_705(c2v_5[70]),
	.c2v_parallelIn_710(c2v_0[71]),
	.c2v_parallelIn_711(c2v_1[71]),
	.c2v_parallelIn_712(c2v_2[71]),
	.c2v_parallelIn_713(c2v_3[71]),
	.c2v_parallelIn_714(c2v_4[71]),
	.c2v_parallelIn_715(c2v_5[71]),
	.c2v_parallelIn_720(c2v_0[72]),
	.c2v_parallelIn_721(c2v_1[72]),
	.c2v_parallelIn_722(c2v_2[72]),
	.c2v_parallelIn_723(c2v_3[72]),
	.c2v_parallelIn_724(c2v_4[72]),
	.c2v_parallelIn_725(c2v_5[72]),
	.c2v_parallelIn_730(c2v_0[73]),
	.c2v_parallelIn_731(c2v_1[73]),
	.c2v_parallelIn_732(c2v_2[73]),
	.c2v_parallelIn_733(c2v_3[73]),
	.c2v_parallelIn_734(c2v_4[73]),
	.c2v_parallelIn_735(c2v_5[73]),
	.c2v_parallelIn_740(c2v_0[74]),
	.c2v_parallelIn_741(c2v_1[74]),
	.c2v_parallelIn_742(c2v_2[74]),
	.c2v_parallelIn_743(c2v_3[74]),
	.c2v_parallelIn_744(c2v_4[74]),
	.c2v_parallelIn_745(c2v_5[74]),
	.c2v_parallelIn_750(c2v_0[75]),
	.c2v_parallelIn_751(c2v_1[75]),
	.c2v_parallelIn_752(c2v_2[75]),
	.c2v_parallelIn_753(c2v_3[75]),
	.c2v_parallelIn_754(c2v_4[75]),
	.c2v_parallelIn_755(c2v_5[75]),
	.c2v_parallelIn_760(c2v_0[76]),
	.c2v_parallelIn_761(c2v_1[76]),
	.c2v_parallelIn_762(c2v_2[76]),
	.c2v_parallelIn_763(c2v_3[76]),
	.c2v_parallelIn_764(c2v_4[76]),
	.c2v_parallelIn_765(c2v_5[76]),
	.c2v_parallelIn_770(c2v_0[77]),
	.c2v_parallelIn_771(c2v_1[77]),
	.c2v_parallelIn_772(c2v_2[77]),
	.c2v_parallelIn_773(c2v_3[77]),
	.c2v_parallelIn_774(c2v_4[77]),
	.c2v_parallelIn_775(c2v_5[77]),
	.c2v_parallelIn_780(c2v_0[78]),
	.c2v_parallelIn_781(c2v_1[78]),
	.c2v_parallelIn_782(c2v_2[78]),
	.c2v_parallelIn_783(c2v_3[78]),
	.c2v_parallelIn_784(c2v_4[78]),
	.c2v_parallelIn_785(c2v_5[78]),
	.c2v_parallelIn_790(c2v_0[79]),
	.c2v_parallelIn_791(c2v_1[79]),
	.c2v_parallelIn_792(c2v_2[79]),
	.c2v_parallelIn_793(c2v_3[79]),
	.c2v_parallelIn_794(c2v_4[79]),
	.c2v_parallelIn_795(c2v_5[79]),
	.c2v_parallelIn_800(c2v_0[80]),
	.c2v_parallelIn_801(c2v_1[80]),
	.c2v_parallelIn_802(c2v_2[80]),
	.c2v_parallelIn_803(c2v_3[80]),
	.c2v_parallelIn_804(c2v_4[80]),
	.c2v_parallelIn_805(c2v_5[80]),
	.c2v_parallelIn_810(c2v_0[81]),
	.c2v_parallelIn_811(c2v_1[81]),
	.c2v_parallelIn_812(c2v_2[81]),
	.c2v_parallelIn_813(c2v_3[81]),
	.c2v_parallelIn_814(c2v_4[81]),
	.c2v_parallelIn_815(c2v_5[81]),
	.c2v_parallelIn_820(c2v_0[82]),
	.c2v_parallelIn_821(c2v_1[82]),
	.c2v_parallelIn_822(c2v_2[82]),
	.c2v_parallelIn_823(c2v_3[82]),
	.c2v_parallelIn_824(c2v_4[82]),
	.c2v_parallelIn_825(c2v_5[82]),
	.c2v_parallelIn_830(c2v_0[83]),
	.c2v_parallelIn_831(c2v_1[83]),
	.c2v_parallelIn_832(c2v_2[83]),
	.c2v_parallelIn_833(c2v_3[83]),
	.c2v_parallelIn_834(c2v_4[83]),
	.c2v_parallelIn_835(c2v_5[83]),
	.c2v_parallelIn_840(c2v_0[84]),
	.c2v_parallelIn_841(c2v_1[84]),
	.c2v_parallelIn_842(c2v_2[84]),
	.c2v_parallelIn_843(c2v_3[84]),
	.c2v_parallelIn_844(c2v_4[84]),
	.c2v_parallelIn_845(c2v_5[84]),
	.c2v_parallelIn_850(c2v_0[85]),
	.c2v_parallelIn_851(c2v_1[85]),
	.c2v_parallelIn_852(c2v_2[85]),
	.c2v_parallelIn_853(c2v_3[85]),
	.c2v_parallelIn_854(c2v_4[85]),
	.c2v_parallelIn_855(c2v_5[85]),
	.c2v_parallelIn_860(c2v_0[86]),
	.c2v_parallelIn_861(c2v_1[86]),
	.c2v_parallelIn_862(c2v_2[86]),
	.c2v_parallelIn_863(c2v_3[86]),
	.c2v_parallelIn_864(c2v_4[86]),
	.c2v_parallelIn_865(c2v_5[86]),
	.c2v_parallelIn_870(c2v_0[87]),
	.c2v_parallelIn_871(c2v_1[87]),
	.c2v_parallelIn_872(c2v_2[87]),
	.c2v_parallelIn_873(c2v_3[87]),
	.c2v_parallelIn_874(c2v_4[87]),
	.c2v_parallelIn_875(c2v_5[87]),
	.c2v_parallelIn_880(c2v_0[88]),
	.c2v_parallelIn_881(c2v_1[88]),
	.c2v_parallelIn_882(c2v_2[88]),
	.c2v_parallelIn_883(c2v_3[88]),
	.c2v_parallelIn_884(c2v_4[88]),
	.c2v_parallelIn_885(c2v_5[88]),
	.c2v_parallelIn_890(c2v_0[89]),
	.c2v_parallelIn_891(c2v_1[89]),
	.c2v_parallelIn_892(c2v_2[89]),
	.c2v_parallelIn_893(c2v_3[89]),
	.c2v_parallelIn_894(c2v_4[89]),
	.c2v_parallelIn_895(c2v_5[89]),
	.c2v_parallelIn_900(c2v_0[90]),
	.c2v_parallelIn_901(c2v_1[90]),
	.c2v_parallelIn_902(c2v_2[90]),
	.c2v_parallelIn_903(c2v_3[90]),
	.c2v_parallelIn_904(c2v_4[90]),
	.c2v_parallelIn_905(c2v_5[90]),
	.c2v_parallelIn_910(c2v_0[91]),
	.c2v_parallelIn_911(c2v_1[91]),
	.c2v_parallelIn_912(c2v_2[91]),
	.c2v_parallelIn_913(c2v_3[91]),
	.c2v_parallelIn_914(c2v_4[91]),
	.c2v_parallelIn_915(c2v_5[91]),
	.c2v_parallelIn_920(c2v_0[92]),
	.c2v_parallelIn_921(c2v_1[92]),
	.c2v_parallelIn_922(c2v_2[92]),
	.c2v_parallelIn_923(c2v_3[92]),
	.c2v_parallelIn_924(c2v_4[92]),
	.c2v_parallelIn_925(c2v_5[92]),
	.c2v_parallelIn_930(c2v_0[93]),
	.c2v_parallelIn_931(c2v_1[93]),
	.c2v_parallelIn_932(c2v_2[93]),
	.c2v_parallelIn_933(c2v_3[93]),
	.c2v_parallelIn_934(c2v_4[93]),
	.c2v_parallelIn_935(c2v_5[93]),
	.c2v_parallelIn_940(c2v_0[94]),
	.c2v_parallelIn_941(c2v_1[94]),
	.c2v_parallelIn_942(c2v_2[94]),
	.c2v_parallelIn_943(c2v_3[94]),
	.c2v_parallelIn_944(c2v_4[94]),
	.c2v_parallelIn_945(c2v_5[94]),
	.c2v_parallelIn_950(c2v_0[95]),
	.c2v_parallelIn_951(c2v_1[95]),
	.c2v_parallelIn_952(c2v_2[95]),
	.c2v_parallelIn_953(c2v_3[95]),
	.c2v_parallelIn_954(c2v_4[95]),
	.c2v_parallelIn_955(c2v_5[95]),
	.c2v_parallelIn_960(c2v_0[96]),
	.c2v_parallelIn_961(c2v_1[96]),
	.c2v_parallelIn_962(c2v_2[96]),
	.c2v_parallelIn_963(c2v_3[96]),
	.c2v_parallelIn_964(c2v_4[96]),
	.c2v_parallelIn_965(c2v_5[96]),
	.c2v_parallelIn_970(c2v_0[97]),
	.c2v_parallelIn_971(c2v_1[97]),
	.c2v_parallelIn_972(c2v_2[97]),
	.c2v_parallelIn_973(c2v_3[97]),
	.c2v_parallelIn_974(c2v_4[97]),
	.c2v_parallelIn_975(c2v_5[97]),
	.c2v_parallelIn_980(c2v_0[98]),
	.c2v_parallelIn_981(c2v_1[98]),
	.c2v_parallelIn_982(c2v_2[98]),
	.c2v_parallelIn_983(c2v_3[98]),
	.c2v_parallelIn_984(c2v_4[98]),
	.c2v_parallelIn_985(c2v_5[98]),
	.c2v_parallelIn_990(c2v_0[99]),
	.c2v_parallelIn_991(c2v_1[99]),
	.c2v_parallelIn_992(c2v_2[99]),
	.c2v_parallelIn_993(c2v_3[99]),
	.c2v_parallelIn_994(c2v_4[99]),
	.c2v_parallelIn_995(c2v_5[99]),
	.c2v_parallelIn_1000(c2v_0[100]),
	.c2v_parallelIn_1001(c2v_1[100]),
	.c2v_parallelIn_1002(c2v_2[100]),
	.c2v_parallelIn_1003(c2v_3[100]),
	.c2v_parallelIn_1004(c2v_4[100]),
	.c2v_parallelIn_1005(c2v_5[100]),
	.c2v_parallelIn_1010(c2v_0[101]),
	.c2v_parallelIn_1011(c2v_1[101]),
	.c2v_parallelIn_1012(c2v_2[101]),
	.c2v_parallelIn_1013(c2v_3[101]),
	.c2v_parallelIn_1014(c2v_4[101]),
	.c2v_parallelIn_1015(c2v_5[101]),
	
	.v2c_parallelIn_00(v2c_0[0]),
	.v2c_parallelIn_01(v2c_1[0]),
	.v2c_parallelIn_02(v2c_2[0]),
	.v2c_parallelIn_10(v2c_0[1]),
	.v2c_parallelIn_11(v2c_1[1]),
	.v2c_parallelIn_12(v2c_2[1]),
	.v2c_parallelIn_20(v2c_0[2]),
	.v2c_parallelIn_21(v2c_1[2]),
	.v2c_parallelIn_22(v2c_2[2]),
	.v2c_parallelIn_30(v2c_0[3]),
	.v2c_parallelIn_31(v2c_1[3]),
	.v2c_parallelIn_32(v2c_2[3]),
	.v2c_parallelIn_40(v2c_0[4]),
	.v2c_parallelIn_41(v2c_1[4]),
	.v2c_parallelIn_42(v2c_2[4]),
	.v2c_parallelIn_50(v2c_0[5]),
	.v2c_parallelIn_51(v2c_1[5]),
	.v2c_parallelIn_52(v2c_2[5]),
	.v2c_parallelIn_60(v2c_0[6]),
	.v2c_parallelIn_61(v2c_1[6]),
	.v2c_parallelIn_62(v2c_2[6]),
	.v2c_parallelIn_70(v2c_0[7]),
	.v2c_parallelIn_71(v2c_1[7]),
	.v2c_parallelIn_72(v2c_2[7]),
	.v2c_parallelIn_80(v2c_0[8]),
	.v2c_parallelIn_81(v2c_1[8]),
	.v2c_parallelIn_82(v2c_2[8]),
	.v2c_parallelIn_90(v2c_0[9]),
	.v2c_parallelIn_91(v2c_1[9]),
	.v2c_parallelIn_92(v2c_2[9]),
	.v2c_parallelIn_100(v2c_0[10]),
	.v2c_parallelIn_101(v2c_1[10]),
	.v2c_parallelIn_102(v2c_2[10]),
	.v2c_parallelIn_110(v2c_0[11]),
	.v2c_parallelIn_111(v2c_1[11]),
	.v2c_parallelIn_112(v2c_2[11]),
	.v2c_parallelIn_120(v2c_0[12]),
	.v2c_parallelIn_121(v2c_1[12]),
	.v2c_parallelIn_122(v2c_2[12]),
	.v2c_parallelIn_130(v2c_0[13]),
	.v2c_parallelIn_131(v2c_1[13]),
	.v2c_parallelIn_132(v2c_2[13]),
	.v2c_parallelIn_140(v2c_0[14]),
	.v2c_parallelIn_141(v2c_1[14]),
	.v2c_parallelIn_142(v2c_2[14]),
	.v2c_parallelIn_150(v2c_0[15]),
	.v2c_parallelIn_151(v2c_1[15]),
	.v2c_parallelIn_152(v2c_2[15]),
	.v2c_parallelIn_160(v2c_0[16]),
	.v2c_parallelIn_161(v2c_1[16]),
	.v2c_parallelIn_162(v2c_2[16]),
	.v2c_parallelIn_170(v2c_0[17]),
	.v2c_parallelIn_171(v2c_1[17]),
	.v2c_parallelIn_172(v2c_2[17]),
	.v2c_parallelIn_180(v2c_0[18]),
	.v2c_parallelIn_181(v2c_1[18]),
	.v2c_parallelIn_182(v2c_2[18]),
	.v2c_parallelIn_190(v2c_0[19]),
	.v2c_parallelIn_191(v2c_1[19]),
	.v2c_parallelIn_192(v2c_2[19]),
	.v2c_parallelIn_200(v2c_0[20]),
	.v2c_parallelIn_201(v2c_1[20]),
	.v2c_parallelIn_202(v2c_2[20]),
	.v2c_parallelIn_210(v2c_0[21]),
	.v2c_parallelIn_211(v2c_1[21]),
	.v2c_parallelIn_212(v2c_2[21]),
	.v2c_parallelIn_220(v2c_0[22]),
	.v2c_parallelIn_221(v2c_1[22]),
	.v2c_parallelIn_222(v2c_2[22]),
	.v2c_parallelIn_230(v2c_0[23]),
	.v2c_parallelIn_231(v2c_1[23]),
	.v2c_parallelIn_232(v2c_2[23]),
	.v2c_parallelIn_240(v2c_0[24]),
	.v2c_parallelIn_241(v2c_1[24]),
	.v2c_parallelIn_242(v2c_2[24]),
	.v2c_parallelIn_250(v2c_0[25]),
	.v2c_parallelIn_251(v2c_1[25]),
	.v2c_parallelIn_252(v2c_2[25]),
	.v2c_parallelIn_260(v2c_0[26]),
	.v2c_parallelIn_261(v2c_1[26]),
	.v2c_parallelIn_262(v2c_2[26]),
	.v2c_parallelIn_270(v2c_0[27]),
	.v2c_parallelIn_271(v2c_1[27]),
	.v2c_parallelIn_272(v2c_2[27]),
	.v2c_parallelIn_280(v2c_0[28]),
	.v2c_parallelIn_281(v2c_1[28]),
	.v2c_parallelIn_282(v2c_2[28]),
	.v2c_parallelIn_290(v2c_0[29]),
	.v2c_parallelIn_291(v2c_1[29]),
	.v2c_parallelIn_292(v2c_2[29]),
	.v2c_parallelIn_300(v2c_0[30]),
	.v2c_parallelIn_301(v2c_1[30]),
	.v2c_parallelIn_302(v2c_2[30]),
	.v2c_parallelIn_310(v2c_0[31]),
	.v2c_parallelIn_311(v2c_1[31]),
	.v2c_parallelIn_312(v2c_2[31]),
	.v2c_parallelIn_320(v2c_0[32]),
	.v2c_parallelIn_321(v2c_1[32]),
	.v2c_parallelIn_322(v2c_2[32]),
	.v2c_parallelIn_330(v2c_0[33]),
	.v2c_parallelIn_331(v2c_1[33]),
	.v2c_parallelIn_332(v2c_2[33]),
	.v2c_parallelIn_340(v2c_0[34]),
	.v2c_parallelIn_341(v2c_1[34]),
	.v2c_parallelIn_342(v2c_2[34]),
	.v2c_parallelIn_350(v2c_0[35]),
	.v2c_parallelIn_351(v2c_1[35]),
	.v2c_parallelIn_352(v2c_2[35]),
	.v2c_parallelIn_360(v2c_0[36]),
	.v2c_parallelIn_361(v2c_1[36]),
	.v2c_parallelIn_362(v2c_2[36]),
	.v2c_parallelIn_370(v2c_0[37]),
	.v2c_parallelIn_371(v2c_1[37]),
	.v2c_parallelIn_372(v2c_2[37]),
	.v2c_parallelIn_380(v2c_0[38]),
	.v2c_parallelIn_381(v2c_1[38]),
	.v2c_parallelIn_382(v2c_2[38]),
	.v2c_parallelIn_390(v2c_0[39]),
	.v2c_parallelIn_391(v2c_1[39]),
	.v2c_parallelIn_392(v2c_2[39]),
	.v2c_parallelIn_400(v2c_0[40]),
	.v2c_parallelIn_401(v2c_1[40]),
	.v2c_parallelIn_402(v2c_2[40]),
	.v2c_parallelIn_410(v2c_0[41]),
	.v2c_parallelIn_411(v2c_1[41]),
	.v2c_parallelIn_412(v2c_2[41]),
	.v2c_parallelIn_420(v2c_0[42]),
	.v2c_parallelIn_421(v2c_1[42]),
	.v2c_parallelIn_422(v2c_2[42]),
	.v2c_parallelIn_430(v2c_0[43]),
	.v2c_parallelIn_431(v2c_1[43]),
	.v2c_parallelIn_432(v2c_2[43]),
	.v2c_parallelIn_440(v2c_0[44]),
	.v2c_parallelIn_441(v2c_1[44]),
	.v2c_parallelIn_442(v2c_2[44]),
	.v2c_parallelIn_450(v2c_0[45]),
	.v2c_parallelIn_451(v2c_1[45]),
	.v2c_parallelIn_452(v2c_2[45]),
	.v2c_parallelIn_460(v2c_0[46]),
	.v2c_parallelIn_461(v2c_1[46]),
	.v2c_parallelIn_462(v2c_2[46]),
	.v2c_parallelIn_470(v2c_0[47]),
	.v2c_parallelIn_471(v2c_1[47]),
	.v2c_parallelIn_472(v2c_2[47]),
	.v2c_parallelIn_480(v2c_0[48]),
	.v2c_parallelIn_481(v2c_1[48]),
	.v2c_parallelIn_482(v2c_2[48]),
	.v2c_parallelIn_490(v2c_0[49]),
	.v2c_parallelIn_491(v2c_1[49]),
	.v2c_parallelIn_492(v2c_2[49]),
	.v2c_parallelIn_500(v2c_0[50]),
	.v2c_parallelIn_501(v2c_1[50]),
	.v2c_parallelIn_502(v2c_2[50]),
	.v2c_parallelIn_510(v2c_0[51]),
	.v2c_parallelIn_511(v2c_1[51]),
	.v2c_parallelIn_512(v2c_2[51]),
	.v2c_parallelIn_520(v2c_0[52]),
	.v2c_parallelIn_521(v2c_1[52]),
	.v2c_parallelIn_522(v2c_2[52]),
	.v2c_parallelIn_530(v2c_0[53]),
	.v2c_parallelIn_531(v2c_1[53]),
	.v2c_parallelIn_532(v2c_2[53]),
	.v2c_parallelIn_540(v2c_0[54]),
	.v2c_parallelIn_541(v2c_1[54]),
	.v2c_parallelIn_542(v2c_2[54]),
	.v2c_parallelIn_550(v2c_0[55]),
	.v2c_parallelIn_551(v2c_1[55]),
	.v2c_parallelIn_552(v2c_2[55]),
	.v2c_parallelIn_560(v2c_0[56]),
	.v2c_parallelIn_561(v2c_1[56]),
	.v2c_parallelIn_562(v2c_2[56]),
	.v2c_parallelIn_570(v2c_0[57]),
	.v2c_parallelIn_571(v2c_1[57]),
	.v2c_parallelIn_572(v2c_2[57]),
	.v2c_parallelIn_580(v2c_0[58]),
	.v2c_parallelIn_581(v2c_1[58]),
	.v2c_parallelIn_582(v2c_2[58]),
	.v2c_parallelIn_590(v2c_0[59]),
	.v2c_parallelIn_591(v2c_1[59]),
	.v2c_parallelIn_592(v2c_2[59]),
	.v2c_parallelIn_600(v2c_0[60]),
	.v2c_parallelIn_601(v2c_1[60]),
	.v2c_parallelIn_602(v2c_2[60]),
	.v2c_parallelIn_610(v2c_0[61]),
	.v2c_parallelIn_611(v2c_1[61]),
	.v2c_parallelIn_612(v2c_2[61]),
	.v2c_parallelIn_620(v2c_0[62]),
	.v2c_parallelIn_621(v2c_1[62]),
	.v2c_parallelIn_622(v2c_2[62]),
	.v2c_parallelIn_630(v2c_0[63]),
	.v2c_parallelIn_631(v2c_1[63]),
	.v2c_parallelIn_632(v2c_2[63]),
	.v2c_parallelIn_640(v2c_0[64]),
	.v2c_parallelIn_641(v2c_1[64]),
	.v2c_parallelIn_642(v2c_2[64]),
	.v2c_parallelIn_650(v2c_0[65]),
	.v2c_parallelIn_651(v2c_1[65]),
	.v2c_parallelIn_652(v2c_2[65]),
	.v2c_parallelIn_660(v2c_0[66]),
	.v2c_parallelIn_661(v2c_1[66]),
	.v2c_parallelIn_662(v2c_2[66]),
	.v2c_parallelIn_670(v2c_0[67]),
	.v2c_parallelIn_671(v2c_1[67]),
	.v2c_parallelIn_672(v2c_2[67]),
	.v2c_parallelIn_680(v2c_0[68]),
	.v2c_parallelIn_681(v2c_1[68]),
	.v2c_parallelIn_682(v2c_2[68]),
	.v2c_parallelIn_690(v2c_0[69]),
	.v2c_parallelIn_691(v2c_1[69]),
	.v2c_parallelIn_692(v2c_2[69]),
	.v2c_parallelIn_700(v2c_0[70]),
	.v2c_parallelIn_701(v2c_1[70]),
	.v2c_parallelIn_702(v2c_2[70]),
	.v2c_parallelIn_710(v2c_0[71]),
	.v2c_parallelIn_711(v2c_1[71]),
	.v2c_parallelIn_712(v2c_2[71]),
	.v2c_parallelIn_720(v2c_0[72]),
	.v2c_parallelIn_721(v2c_1[72]),
	.v2c_parallelIn_722(v2c_2[72]),
	.v2c_parallelIn_730(v2c_0[73]),
	.v2c_parallelIn_731(v2c_1[73]),
	.v2c_parallelIn_732(v2c_2[73]),
	.v2c_parallelIn_740(v2c_0[74]),
	.v2c_parallelIn_741(v2c_1[74]),
	.v2c_parallelIn_742(v2c_2[74]),
	.v2c_parallelIn_750(v2c_0[75]),
	.v2c_parallelIn_751(v2c_1[75]),
	.v2c_parallelIn_752(v2c_2[75]),
	.v2c_parallelIn_760(v2c_0[76]),
	.v2c_parallelIn_761(v2c_1[76]),
	.v2c_parallelIn_762(v2c_2[76]),
	.v2c_parallelIn_770(v2c_0[77]),
	.v2c_parallelIn_771(v2c_1[77]),
	.v2c_parallelIn_772(v2c_2[77]),
	.v2c_parallelIn_780(v2c_0[78]),
	.v2c_parallelIn_781(v2c_1[78]),
	.v2c_parallelIn_782(v2c_2[78]),
	.v2c_parallelIn_790(v2c_0[79]),
	.v2c_parallelIn_791(v2c_1[79]),
	.v2c_parallelIn_792(v2c_2[79]),
	.v2c_parallelIn_800(v2c_0[80]),
	.v2c_parallelIn_801(v2c_1[80]),
	.v2c_parallelIn_802(v2c_2[80]),
	.v2c_parallelIn_810(v2c_0[81]),
	.v2c_parallelIn_811(v2c_1[81]),
	.v2c_parallelIn_812(v2c_2[81]),
	.v2c_parallelIn_820(v2c_0[82]),
	.v2c_parallelIn_821(v2c_1[82]),
	.v2c_parallelIn_822(v2c_2[82]),
	.v2c_parallelIn_830(v2c_0[83]),
	.v2c_parallelIn_831(v2c_1[83]),
	.v2c_parallelIn_832(v2c_2[83]),
	.v2c_parallelIn_840(v2c_0[84]),
	.v2c_parallelIn_841(v2c_1[84]),
	.v2c_parallelIn_842(v2c_2[84]),
	.v2c_parallelIn_850(v2c_0[85]),
	.v2c_parallelIn_851(v2c_1[85]),
	.v2c_parallelIn_852(v2c_2[85]),
	.v2c_parallelIn_860(v2c_0[86]),
	.v2c_parallelIn_861(v2c_1[86]),
	.v2c_parallelIn_862(v2c_2[86]),
	.v2c_parallelIn_870(v2c_0[87]),
	.v2c_parallelIn_871(v2c_1[87]),
	.v2c_parallelIn_872(v2c_2[87]),
	.v2c_parallelIn_880(v2c_0[88]),
	.v2c_parallelIn_881(v2c_1[88]),
	.v2c_parallelIn_882(v2c_2[88]),
	.v2c_parallelIn_890(v2c_0[89]),
	.v2c_parallelIn_891(v2c_1[89]),
	.v2c_parallelIn_892(v2c_2[89]),
	.v2c_parallelIn_900(v2c_0[90]),
	.v2c_parallelIn_901(v2c_1[90]),
	.v2c_parallelIn_902(v2c_2[90]),
	.v2c_parallelIn_910(v2c_0[91]),
	.v2c_parallelIn_911(v2c_1[91]),
	.v2c_parallelIn_912(v2c_2[91]),
	.v2c_parallelIn_920(v2c_0[92]),
	.v2c_parallelIn_921(v2c_1[92]),
	.v2c_parallelIn_922(v2c_2[92]),
	.v2c_parallelIn_930(v2c_0[93]),
	.v2c_parallelIn_931(v2c_1[93]),
	.v2c_parallelIn_932(v2c_2[93]),
	.v2c_parallelIn_940(v2c_0[94]),
	.v2c_parallelIn_941(v2c_1[94]),
	.v2c_parallelIn_942(v2c_2[94]),
	.v2c_parallelIn_950(v2c_0[95]),
	.v2c_parallelIn_951(v2c_1[95]),
	.v2c_parallelIn_952(v2c_2[95]),
	.v2c_parallelIn_960(v2c_0[96]),
	.v2c_parallelIn_961(v2c_1[96]),
	.v2c_parallelIn_962(v2c_2[96]),
	.v2c_parallelIn_970(v2c_0[97]),
	.v2c_parallelIn_971(v2c_1[97]),
	.v2c_parallelIn_972(v2c_2[97]),
	.v2c_parallelIn_980(v2c_0[98]),
	.v2c_parallelIn_981(v2c_1[98]),
	.v2c_parallelIn_982(v2c_2[98]),
	.v2c_parallelIn_990(v2c_0[99]),
	.v2c_parallelIn_991(v2c_1[99]),
	.v2c_parallelIn_992(v2c_2[99]),
	.v2c_parallelIn_1000(v2c_0[100]),
	.v2c_parallelIn_1001(v2c_1[100]),
	.v2c_parallelIn_1002(v2c_2[100]),
	.v2c_parallelIn_1010(v2c_0[101]),
	.v2c_parallelIn_1011(v2c_1[101]),
	.v2c_parallelIn_1012(v2c_2[101]),
	.v2c_parallelIn_1020(v2c_0[102]),
	.v2c_parallelIn_1021(v2c_1[102]),
	.v2c_parallelIn_1022(v2c_2[102]),
	.v2c_parallelIn_1030(v2c_0[103]),
	.v2c_parallelIn_1031(v2c_1[103]),
	.v2c_parallelIn_1032(v2c_2[103]),
	.v2c_parallelIn_1040(v2c_0[104]),
	.v2c_parallelIn_1041(v2c_1[104]),
	.v2c_parallelIn_1042(v2c_2[104]),
	.v2c_parallelIn_1050(v2c_0[105]),
	.v2c_parallelIn_1051(v2c_1[105]),
	.v2c_parallelIn_1052(v2c_2[105]),
	.v2c_parallelIn_1060(v2c_0[106]),
	.v2c_parallelIn_1061(v2c_1[106]),
	.v2c_parallelIn_1062(v2c_2[106]),
	.v2c_parallelIn_1070(v2c_0[107]),
	.v2c_parallelIn_1071(v2c_1[107]),
	.v2c_parallelIn_1072(v2c_2[107]),
	.v2c_parallelIn_1080(v2c_0[108]),
	.v2c_parallelIn_1081(v2c_1[108]),
	.v2c_parallelIn_1082(v2c_2[108]),
	.v2c_parallelIn_1090(v2c_0[109]),
	.v2c_parallelIn_1091(v2c_1[109]),
	.v2c_parallelIn_1092(v2c_2[109]),
	.v2c_parallelIn_1100(v2c_0[110]),
	.v2c_parallelIn_1101(v2c_1[110]),
	.v2c_parallelIn_1102(v2c_2[110]),
	.v2c_parallelIn_1110(v2c_0[111]),
	.v2c_parallelIn_1111(v2c_1[111]),
	.v2c_parallelIn_1112(v2c_2[111]),
	.v2c_parallelIn_1120(v2c_0[112]),
	.v2c_parallelIn_1121(v2c_1[112]),
	.v2c_parallelIn_1122(v2c_2[112]),
	.v2c_parallelIn_1130(v2c_0[113]),
	.v2c_parallelIn_1131(v2c_1[113]),
	.v2c_parallelIn_1132(v2c_2[113]),
	.v2c_parallelIn_1140(v2c_0[114]),
	.v2c_parallelIn_1141(v2c_1[114]),
	.v2c_parallelIn_1142(v2c_2[114]),
	.v2c_parallelIn_1150(v2c_0[115]),
	.v2c_parallelIn_1151(v2c_1[115]),
	.v2c_parallelIn_1152(v2c_2[115]),
	.v2c_parallelIn_1160(v2c_0[116]),
	.v2c_parallelIn_1161(v2c_1[116]),
	.v2c_parallelIn_1162(v2c_2[116]),
	.v2c_parallelIn_1170(v2c_0[117]),
	.v2c_parallelIn_1171(v2c_1[117]),
	.v2c_parallelIn_1172(v2c_2[117]),
	.v2c_parallelIn_1180(v2c_0[118]),
	.v2c_parallelIn_1181(v2c_1[118]),
	.v2c_parallelIn_1182(v2c_2[118]),
	.v2c_parallelIn_1190(v2c_0[119]),
	.v2c_parallelIn_1191(v2c_1[119]),
	.v2c_parallelIn_1192(v2c_2[119]),
	.v2c_parallelIn_1200(v2c_0[120]),
	.v2c_parallelIn_1201(v2c_1[120]),
	.v2c_parallelIn_1202(v2c_2[120]),
	.v2c_parallelIn_1210(v2c_0[121]),
	.v2c_parallelIn_1211(v2c_1[121]),
	.v2c_parallelIn_1212(v2c_2[121]),
	.v2c_parallelIn_1220(v2c_0[122]),
	.v2c_parallelIn_1221(v2c_1[122]),
	.v2c_parallelIn_1222(v2c_2[122]),
	.v2c_parallelIn_1230(v2c_0[123]),
	.v2c_parallelIn_1231(v2c_1[123]),
	.v2c_parallelIn_1232(v2c_2[123]),
	.v2c_parallelIn_1240(v2c_0[124]),
	.v2c_parallelIn_1241(v2c_1[124]),
	.v2c_parallelIn_1242(v2c_2[124]),
	.v2c_parallelIn_1250(v2c_0[125]),
	.v2c_parallelIn_1251(v2c_1[125]),
	.v2c_parallelIn_1252(v2c_2[125]),
	.v2c_parallelIn_1260(v2c_0[126]),
	.v2c_parallelIn_1261(v2c_1[126]),
	.v2c_parallelIn_1262(v2c_2[126]),
	.v2c_parallelIn_1270(v2c_0[127]),
	.v2c_parallelIn_1271(v2c_1[127]),
	.v2c_parallelIn_1272(v2c_2[127]),
	.v2c_parallelIn_1280(v2c_0[128]),
	.v2c_parallelIn_1281(v2c_1[128]),
	.v2c_parallelIn_1282(v2c_2[128]),
	.v2c_parallelIn_1290(v2c_0[129]),
	.v2c_parallelIn_1291(v2c_1[129]),
	.v2c_parallelIn_1292(v2c_2[129]),
	.v2c_parallelIn_1300(v2c_0[130]),
	.v2c_parallelIn_1301(v2c_1[130]),
	.v2c_parallelIn_1302(v2c_2[130]),
	.v2c_parallelIn_1310(v2c_0[131]),
	.v2c_parallelIn_1311(v2c_1[131]),
	.v2c_parallelIn_1312(v2c_2[131]),
	.v2c_parallelIn_1320(v2c_0[132]),
	.v2c_parallelIn_1321(v2c_1[132]),
	.v2c_parallelIn_1322(v2c_2[132]),
	.v2c_parallelIn_1330(v2c_0[133]),
	.v2c_parallelIn_1331(v2c_1[133]),
	.v2c_parallelIn_1332(v2c_2[133]),
	.v2c_parallelIn_1340(v2c_0[134]),
	.v2c_parallelIn_1341(v2c_1[134]),
	.v2c_parallelIn_1342(v2c_2[134]),
	.v2c_parallelIn_1350(v2c_0[135]),
	.v2c_parallelIn_1351(v2c_1[135]),
	.v2c_parallelIn_1352(v2c_2[135]),
	.v2c_parallelIn_1360(v2c_0[136]),
	.v2c_parallelIn_1361(v2c_1[136]),
	.v2c_parallelIn_1362(v2c_2[136]),
	.v2c_parallelIn_1370(v2c_0[137]),
	.v2c_parallelIn_1371(v2c_1[137]),
	.v2c_parallelIn_1372(v2c_2[137]),
	.v2c_parallelIn_1380(v2c_0[138]),
	.v2c_parallelIn_1381(v2c_1[138]),
	.v2c_parallelIn_1382(v2c_2[138]),
	.v2c_parallelIn_1390(v2c_0[139]),
	.v2c_parallelIn_1391(v2c_1[139]),
	.v2c_parallelIn_1392(v2c_2[139]),
	.v2c_parallelIn_1400(v2c_0[140]),
	.v2c_parallelIn_1401(v2c_1[140]),
	.v2c_parallelIn_1402(v2c_2[140]),
	.v2c_parallelIn_1410(v2c_0[141]),
	.v2c_parallelIn_1411(v2c_1[141]),
	.v2c_parallelIn_1412(v2c_2[141]),
	.v2c_parallelIn_1420(v2c_0[142]),
	.v2c_parallelIn_1421(v2c_1[142]),
	.v2c_parallelIn_1422(v2c_2[142]),
	.v2c_parallelIn_1430(v2c_0[143]),
	.v2c_parallelIn_1431(v2c_1[143]),
	.v2c_parallelIn_1432(v2c_2[143]),
	.v2c_parallelIn_1440(v2c_0[144]),
	.v2c_parallelIn_1441(v2c_1[144]),
	.v2c_parallelIn_1442(v2c_2[144]),
	.v2c_parallelIn_1450(v2c_0[145]),
	.v2c_parallelIn_1451(v2c_1[145]),
	.v2c_parallelIn_1452(v2c_2[145]),
	.v2c_parallelIn_1460(v2c_0[146]),
	.v2c_parallelIn_1461(v2c_1[146]),
	.v2c_parallelIn_1462(v2c_2[146]),
	.v2c_parallelIn_1470(v2c_0[147]),
	.v2c_parallelIn_1471(v2c_1[147]),
	.v2c_parallelIn_1472(v2c_2[147]),
	.v2c_parallelIn_1480(v2c_0[148]),
	.v2c_parallelIn_1481(v2c_1[148]),
	.v2c_parallelIn_1482(v2c_2[148]),
	.v2c_parallelIn_1490(v2c_0[149]),
	.v2c_parallelIn_1491(v2c_1[149]),
	.v2c_parallelIn_1492(v2c_2[149]),
	.v2c_parallelIn_1500(v2c_0[150]),
	.v2c_parallelIn_1501(v2c_1[150]),
	.v2c_parallelIn_1502(v2c_2[150]),
	.v2c_parallelIn_1510(v2c_0[151]),
	.v2c_parallelIn_1511(v2c_1[151]),
	.v2c_parallelIn_1512(v2c_2[151]),
	.v2c_parallelIn_1520(v2c_0[152]),
	.v2c_parallelIn_1521(v2c_1[152]),
	.v2c_parallelIn_1522(v2c_2[152]),
	.v2c_parallelIn_1530(v2c_0[153]),
	.v2c_parallelIn_1531(v2c_1[153]),
	.v2c_parallelIn_1532(v2c_2[153]),
	.v2c_parallelIn_1540(v2c_0[154]),
	.v2c_parallelIn_1541(v2c_1[154]),
	.v2c_parallelIn_1542(v2c_2[154]),
	.v2c_parallelIn_1550(v2c_0[155]),
	.v2c_parallelIn_1551(v2c_1[155]),
	.v2c_parallelIn_1552(v2c_2[155]),
	.v2c_parallelIn_1560(v2c_0[156]),
	.v2c_parallelIn_1561(v2c_1[156]),
	.v2c_parallelIn_1562(v2c_2[156]),
	.v2c_parallelIn_1570(v2c_0[157]),
	.v2c_parallelIn_1571(v2c_1[157]),
	.v2c_parallelIn_1572(v2c_2[157]),
	.v2c_parallelIn_1580(v2c_0[158]),
	.v2c_parallelIn_1581(v2c_1[158]),
	.v2c_parallelIn_1582(v2c_2[158]),
	.v2c_parallelIn_1590(v2c_0[159]),
	.v2c_parallelIn_1591(v2c_1[159]),
	.v2c_parallelIn_1592(v2c_2[159]),
	.v2c_parallelIn_1600(v2c_0[160]),
	.v2c_parallelIn_1601(v2c_1[160]),
	.v2c_parallelIn_1602(v2c_2[160]),
	.v2c_parallelIn_1610(v2c_0[161]),
	.v2c_parallelIn_1611(v2c_1[161]),
	.v2c_parallelIn_1612(v2c_2[161]),
	.v2c_parallelIn_1620(v2c_0[162]),
	.v2c_parallelIn_1621(v2c_1[162]),
	.v2c_parallelIn_1622(v2c_2[162]),
	.v2c_parallelIn_1630(v2c_0[163]),
	.v2c_parallelIn_1631(v2c_1[163]),
	.v2c_parallelIn_1632(v2c_2[163]),
	.v2c_parallelIn_1640(v2c_0[164]),
	.v2c_parallelIn_1641(v2c_1[164]),
	.v2c_parallelIn_1642(v2c_2[164]),
	.v2c_parallelIn_1650(v2c_0[165]),
	.v2c_parallelIn_1651(v2c_1[165]),
	.v2c_parallelIn_1652(v2c_2[165]),
	.v2c_parallelIn_1660(v2c_0[166]),
	.v2c_parallelIn_1661(v2c_1[166]),
	.v2c_parallelIn_1662(v2c_2[166]),
	.v2c_parallelIn_1670(v2c_0[167]),
	.v2c_parallelIn_1671(v2c_1[167]),
	.v2c_parallelIn_1672(v2c_2[167]),
	.v2c_parallelIn_1680(v2c_0[168]),
	.v2c_parallelIn_1681(v2c_1[168]),
	.v2c_parallelIn_1682(v2c_2[168]),
	.v2c_parallelIn_1690(v2c_0[169]),
	.v2c_parallelIn_1691(v2c_1[169]),
	.v2c_parallelIn_1692(v2c_2[169]),
	.v2c_parallelIn_1700(v2c_0[170]),
	.v2c_parallelIn_1701(v2c_1[170]),
	.v2c_parallelIn_1702(v2c_2[170]),
	.v2c_parallelIn_1710(v2c_0[171]),
	.v2c_parallelIn_1711(v2c_1[171]),
	.v2c_parallelIn_1712(v2c_2[171]),
	.v2c_parallelIn_1720(v2c_0[172]),
	.v2c_parallelIn_1721(v2c_1[172]),
	.v2c_parallelIn_1722(v2c_2[172]),
	.v2c_parallelIn_1730(v2c_0[173]),
	.v2c_parallelIn_1731(v2c_1[173]),
	.v2c_parallelIn_1732(v2c_2[173]),
	.v2c_parallelIn_1740(v2c_0[174]),
	.v2c_parallelIn_1741(v2c_1[174]),
	.v2c_parallelIn_1742(v2c_2[174]),
	.v2c_parallelIn_1750(v2c_0[175]),
	.v2c_parallelIn_1751(v2c_1[175]),
	.v2c_parallelIn_1752(v2c_2[175]),
	.v2c_parallelIn_1760(v2c_0[176]),
	.v2c_parallelIn_1761(v2c_1[176]),
	.v2c_parallelIn_1762(v2c_2[176]),
	.v2c_parallelIn_1770(v2c_0[177]),
	.v2c_parallelIn_1771(v2c_1[177]),
	.v2c_parallelIn_1772(v2c_2[177]),
	.v2c_parallelIn_1780(v2c_0[178]),
	.v2c_parallelIn_1781(v2c_1[178]),
	.v2c_parallelIn_1782(v2c_2[178]),
	.v2c_parallelIn_1790(v2c_0[179]),
	.v2c_parallelIn_1791(v2c_1[179]),
	.v2c_parallelIn_1792(v2c_2[179]),
	.v2c_parallelIn_1800(v2c_0[180]),
	.v2c_parallelIn_1801(v2c_1[180]),
	.v2c_parallelIn_1802(v2c_2[180]),
	.v2c_parallelIn_1810(v2c_0[181]),
	.v2c_parallelIn_1811(v2c_1[181]),
	.v2c_parallelIn_1812(v2c_2[181]),
	.v2c_parallelIn_1820(v2c_0[182]),
	.v2c_parallelIn_1821(v2c_1[182]),
	.v2c_parallelIn_1822(v2c_2[182]),
	.v2c_parallelIn_1830(v2c_0[183]),
	.v2c_parallelIn_1831(v2c_1[183]),
	.v2c_parallelIn_1832(v2c_2[183]),
	.v2c_parallelIn_1840(v2c_0[184]),
	.v2c_parallelIn_1841(v2c_1[184]),
	.v2c_parallelIn_1842(v2c_2[184]),
	.v2c_parallelIn_1850(v2c_0[185]),
	.v2c_parallelIn_1851(v2c_1[185]),
	.v2c_parallelIn_1852(v2c_2[185]),
	.v2c_parallelIn_1860(v2c_0[186]),
	.v2c_parallelIn_1861(v2c_1[186]),
	.v2c_parallelIn_1862(v2c_2[186]),
	.v2c_parallelIn_1870(v2c_0[187]),
	.v2c_parallelIn_1871(v2c_1[187]),
	.v2c_parallelIn_1872(v2c_2[187]),
	.v2c_parallelIn_1880(v2c_0[188]),
	.v2c_parallelIn_1881(v2c_1[188]),
	.v2c_parallelIn_1882(v2c_2[188]),
	.v2c_parallelIn_1890(v2c_0[189]),
	.v2c_parallelIn_1891(v2c_1[189]),
	.v2c_parallelIn_1892(v2c_2[189]),
	.v2c_parallelIn_1900(v2c_0[190]),
	.v2c_parallelIn_1901(v2c_1[190]),
	.v2c_parallelIn_1902(v2c_2[190]),
	.v2c_parallelIn_1910(v2c_0[191]),
	.v2c_parallelIn_1911(v2c_1[191]),
	.v2c_parallelIn_1912(v2c_2[191]),
	.v2c_parallelIn_1920(v2c_0[192]),
	.v2c_parallelIn_1921(v2c_1[192]),
	.v2c_parallelIn_1922(v2c_2[192]),
	.v2c_parallelIn_1930(v2c_0[193]),
	.v2c_parallelIn_1931(v2c_1[193]),
	.v2c_parallelIn_1932(v2c_2[193]),
	.v2c_parallelIn_1940(v2c_0[194]),
	.v2c_parallelIn_1941(v2c_1[194]),
	.v2c_parallelIn_1942(v2c_2[194]),
	.v2c_parallelIn_1950(v2c_0[195]),
	.v2c_parallelIn_1951(v2c_1[195]),
	.v2c_parallelIn_1952(v2c_2[195]),
	.v2c_parallelIn_1960(v2c_0[196]),
	.v2c_parallelIn_1961(v2c_1[196]),
	.v2c_parallelIn_1962(v2c_2[196]),
	.v2c_parallelIn_1970(v2c_0[197]),
	.v2c_parallelIn_1971(v2c_1[197]),
	.v2c_parallelIn_1972(v2c_2[197]),
	.v2c_parallelIn_1980(v2c_0[198]),
	.v2c_parallelIn_1981(v2c_1[198]),
	.v2c_parallelIn_1982(v2c_2[198]),
	.v2c_parallelIn_1990(v2c_0[199]),
	.v2c_parallelIn_1991(v2c_1[199]),
	.v2c_parallelIn_1992(v2c_2[199]),
	.v2c_parallelIn_2000(v2c_0[200]),
	.v2c_parallelIn_2001(v2c_1[200]),
	.v2c_parallelIn_2002(v2c_2[200]),
	.v2c_parallelIn_2010(v2c_0[201]),
	.v2c_parallelIn_2011(v2c_1[201]),
	.v2c_parallelIn_2012(v2c_2[201]),
	.v2c_parallelIn_2020(v2c_0[202]),
	.v2c_parallelIn_2021(v2c_1[202]),
	.v2c_parallelIn_2022(v2c_2[202]),
	.v2c_parallelIn_2030(v2c_0[203]),
	.v2c_parallelIn_2031(v2c_1[203]),
	.v2c_parallelIn_2032(v2c_2[203]),
	
	.load({v2c_load[0], c2v_load[0]}),
	.parallel_en ({v2c_msg_en[0], c2v_msg_en[0]}),
	.serial_clk (read_clk)
};

/*
halfDuplex_parallel2serial #(
	.MSG_WIDTH(`DATAPATH_WIDTH) // the default bit widith of one message is 4-bit
) cnu_interface_u0(
    .serial_inout (extrinsic_route),
    .parallel_out (v2c_parallel_out[`DATAPATH_WIDTH-1:0]),
    
    .parallel_in (c2v_parallel_in[`DATAPATH_WIDTH-1:0]),
    .load		 (c2v_load[0]),
    .parallel_en (c2v_msg_en[0]), // to decide the direction of serial_inout port, i.e., '0' -> input whilst '1' -> output
    .sys_clk (read_clk)
);
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) c2v_parallel_in <= 10;
	else if(sys_fsm_state[0] == 4) c2v_parallel_in <= c2v_parallel_in + 1;
end
*/
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) c2v_msg_busy <= 0;
	else c2v_msg_busy <= c2v_msg_en[0];
end
assign c2v_latch_en = {c2v_msg_busy && ~c2v_msg_en[0]}; // the busy sign of PSP: 00b -> idle, 01b -> load, 11b -> message passing, 10b -> message passing finished

always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) 
		c2v_latch[`DATAPATH_WIDTH-1:0] <= 0;
	else if(c2v_latch_en == 1'b1) 
		c2v_latch[`DATAPATH_WIDTH-1:0] <= c2v_parallel_out[`DATAPATH_WIDTH-1:0];
	else 
		c2v_latch[`DATAPATH_WIDTH-1:0] <= c2v_latch[`DATAPATH_WIDTH-1:0];
end
/*
halfDuplex_parallel2serial #(
	.MSG_WIDTH(`DATAPATH_WIDTH) // the default bit widith of one message is 4-bit
) vnu_interface_u0(
    .serial_inout (extrinsic_route),
    .parallel_out (c2v_parallel_out[`DATAPATH_WIDTH-1:0]),
    
    .parallel_in (v2c_parallel_in[`DATAPATH_WIDTH-1:0]),
    .load		 (v2c_load[0]),
    .parallel_en (v2c_msg_en[0]), // to decide the direction of serial_inout port, i.e., '0' -> input whilst '1' -> output
    .sys_clk (read_clk)
);
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) v2c_parallel_in <= 1;
	else if(sys_fsm_state[0] == 8) v2c_parallel_in <= v2c_parallel_in + 1;
end
*/
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) v2c_msg_busy <= 0;
	else v2c_msg_busy <= v2c_msg_en[0];
end
assign v2c_latch_en = {v2c_msg_busy && ~v2c_msg_en[0]}; // the busy sign of PSP: 00b -> idle, 01b -> load, 11b -> message passing, 10b -> message passing finished

always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) 
		v2c_latch[`DATAPATH_WIDTH-1:0] <= 0;
	else if(v2c_latch_en == 1'b1) 
		v2c_latch[`DATAPATH_WIDTH-1:0] <= v2c_parallel_out[`DATAPATH_WIDTH-1:0];
	else 
		v2c_latch[`DATAPATH_WIDTH-1:0] <= v2c_latch[`DATAPATH_WIDTH-1:0];
end
//////////////////////////////////////////////////////////////////////////////////////////////////////
initial begin
       $dumpfile("sys_fsm.vcd");
       $dumpvars;
end

initial begin
	#0 read_clk     <= 1'b0;
	#2.5;
	forever #5   read_clk     <= ~read_clk;
end
initial begin
	#0 cn_write_clk <= 1'b0;
	//#2.5;
	forever #2.5 cn_write_clk <= ~cn_write_clk;
end
initial begin
	#0 vn_write_clk <= 1'b0;
	forever #2.5 vn_write_clk <= ~vn_write_clk;
end
initial begin
	#0 dn_write_clk <= 1'b0;
	forever #2.5 dn_write_clk <= ~dn_write_clk;
end
initial begin
	#0;
	rstn <= 1'b0;
	
	#2.5;
	#(10*100);
	rstn <= 1'b1;
end

/*
reg [3:0] iter_cnt [0:1];
initial #0 iter_cnt[0] <= 4'd0;
always @(posedge read_clk) begin
	if(sys_fsm_state[0] == P2P_V_OUT) iter_cnt[0] <= iter_cnt[0] + 1'b1;
	else if(iter_cnt[0] == 5) iter_cnt[0] <= 4'd0;
end 
initial #0 iter_cnt[1] <= 4'd0;
always @(posedge read_clk) begin
	if(sys_fsm_state[1] == P2P_V_OUT) iter_cnt[1] <= iter_cnt[1] + 1'b1;
	else if(iter_cnt[1] == 5) iter_cnt[1] <= 4'd0;
end 
initial #0 iter_termination[INTER_FRAME_LEVEL-1:0] <= 'd0;
always @(posedge read_clk) begin
	if(iter_cnt[0] == 5 && sys_fsm_state[0] == CNU_PIPE && de_frame_start[0]) iter_termination[0] <= 1'b1;
	else if(de_frame_start[0] == 1'b1 && iter_termination[0] == 1'b1) iter_termination[0] <= 1'b0;  
end
always @(posedge read_clk) begin
	if(iter_cnt[1] == 5 && sys_fsm_state[1] == CNU_PIPE && de_frame_start[1]) iter_termination[1] <= 1'b1;
	else if(de_frame_start[1] == 1'b1 && iter_termination[1] == 1'b1) iter_termination[1] <= 1'b0;  
end
*/

always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) 
		iter_cnt <= 0;
	else if(sys_fsm_state[0] == VNU_OUT)
		iter_cnt <= iter_cnt + 1'b1;
	else if(iter_termination[0] == 1'b1)
		iter_cnt <= 0;
	else
		iter_cnt <= iter_cnt;
end

reg [1:0] termination_latch;
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) termination_latch <= 0;
	else termination_latch[1:0] <= {termination_latch[0], iter_termination[0]};
end
always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) codeword_cnt <= 0;
	else if(termination_latch[1:0] == 2'b01) codeword_cnt <= codeword_cnt + 1'b1;
end

//////////////////////////////////////////////////////////////////////////////////////////////////////
// Log File
//integer fsm_log;
//initial fsm_log = $fopen("fsm_log.txt","w");
//always @(posedge read_clk) begin
//    if(rstn) begin
//		case (sys_fsm_state[0])
//			INIT_LOAD: $fwrite(fsm_log,"INIT_LOAD\t\t");
//			LLR_FETCH: $fwrite(fsm_log,"LLR_FETCH\t");
//			LLR_FETCH_OUT: $fwrite(fsm_log,"LLR_FETCH_OUT\t");
//			CNU_PIPE: $fwrite(fsm_log,"CNU_PIPE\t");
//			CNU_OUT: $fwrite(fsm_log,"CNU_OUT\t\t");
//			P2P_C: $fwrite(fsm_log,"P2P_C\t\t");
//			P2P_C_OUT: $fwrite(fsm_log,"P2P_C_OUT\t");
//			VNU_PIPE: $fwrite(fsm_log,"VNU_PIPE\t");
//			VNU_OUT: $fwrite(fsm_log,"VNU_OUT\t\t");
//			P2P_V: $fwrite(fsm_log,"P2P_V\t\t");
//			P2P_V_OUT: $fwrite(fsm_log,"(Iter%d)P2P_V_OUT\t", iter_cnt[0]);
//		endcase
//		/*
//		case (sys_fsm_state[1])
//			INIT_LOAD: $fwrite(fsm_log,"CONFIG");
//			LLR_FETCH: $fwrite(fsm_log,"LLR_FETCH");
//			LLR_FETCH_OUT: $fwrite(fsm_log,"LLR_FETCH_OUT");
//			CNU_PIPE: $fwrite(fsm_log,"CNU_PIPE");
//			CNU_OUT: $fwrite(fsm_log,"CNU_OUT");
//			P2P_C: $fwrite(fsm_log,"P2P_C");
//			P2P_C_OUT: $fwrite(fsm_log,"P2P_C_OUT");
//			VNU_PIPE: $fwrite(fsm_log,"VNU_PIPE");
//			VNU_OUT: $fwrite(fsm_log,"VNU_OUT");
//			P2P_V: $fwrite(fsm_log,"P2P_V");
//			P2P_V_OUT: $fwrite(fsm_log,"(Iter%d)P2P_V_OUT", iter_cnt[1]);
//		endcase
//		*/
//		$fwrite(fsm_log, "\tcn_we: (%b)\tvn_we: (%b)\tdn_we: (%b)\n", fsm_cn_ram_we[0], fsm_vn_ram_we[0], fsm_dn_ram_we[0]);
//    end 
//end
//
//integer fsm_out [0:1];
//initial begin
//	fsm_out[0] = $fopen("fsm_out.0.txt", "w");
//	fsm_out[1] = $fopen("fsm_out.1.txt", "w");
//end
//always @(posedge read_clk) begin
//	if(rstn) begin
//	    $fwrite(fsm_out[0], "iter_termination:%d, llr_fetch:%d, v2c_src:%d, v2c_msg:%d, cnu_rd:%d, c2v_msg_en:%d, vnu_rd:%d, inter_frame_en:%d, de_frame_start:%d\n", 
//			iter_termination[0], 
//			llr_fetch[0],
//			v2c_src[0],
//			v2c_msg_en[0],
//			cnu_rd[0],
//			c2v_msg_en[0],
//			vnu_rd[0],
//			inter_frame_en[0],
//			de_frame_start[0]
//	    );
//		/*
//	    $fwrite(fsm_out[1], "iter_termination:%d, llr_fetch:%d, v2c_src:%d, v2c_msg:%d, cnu_rd:%d, c2v_msg_en:%d, vnu_rd:%d, inter_frame_en:%d, de_frame_start:%d\n", 
//			iter_termination[1], 
//			llr_fetch[1],
//			v2c_src[1],
//			v2c_msg_en[1],
//			cnu_rd[1],
//			c2v_msg_en[1],
//			vnu_rd[1],
//			inter_frame_en[1],
//			de_frame_start[1]
//	    );
//		*/
//	end
//end
//
//// Log files of write-enable signals for IB-CNU and IB-VNU RAMs
//integer fsm_we_out [0:1];
//initial begin
//	fsm_we_out[0] = $fopen("cnu_we.txt", "w");
//	//fsm_we_out[1] = $fopen("vnu_we.txt", "w");
//end
//always @(posedge read_clk) begin
//	if(rstn) begin
//	    $fwrite(fsm_we_out[0], "(%b, %b)\n", fsm_cn_ram_we[0], fsm_cn_ram_we[1]);
//	    //$fwrite(fsm_we_out[1], "(%b, %b)\n", fsm_vn_ram_we[0], fsm_vn_ram_we[1]);
//	end
//end
//////////////////////////////////////////////////////////////////////////////////////////////////////

always @(posedge read_clk, negedge rstn) begin
	if(rstn == 1'b0) iter_termination <= 0;
	else if(iter_cnt == simulate_iteration) iter_termination <= 2'b11;
	else if(iter_termination == 2'b11) iter_termination <= 0;
end

initial begin
	wait(codeword_cnt == simulate_codewords);  //#(10*144);
	#20;
	//#500000;

	//$fclose(fsm_log);
	//$fclose(fsm_out[0]);
	////$fclose(fsm_out[1]);
	//$fclose(fsm_we_out[0]);
	////$fclose(fsm_we_out[1]);
    $finish;
end
endmodule
