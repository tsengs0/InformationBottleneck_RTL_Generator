`include "define.vh"

`ifdef SCHED_4_6
module ram_pageAlign_interface_submatrix_4#(
	parameter QUAN_SIZE = 4,
	parameter CHECK_PARALLELISM = 255,
	parameter LAYER_NUM = 3
) (
	output wire [QUAN_SIZE-1:0] msg_out_0,
	output wire [QUAN_SIZE-1:0] msg_out_1,
	output wire [QUAN_SIZE-1:0] msg_out_2,
	output wire [QUAN_SIZE-1:0] msg_out_3,
	output wire [QUAN_SIZE-1:0] msg_out_4,
	output wire [QUAN_SIZE-1:0] msg_out_5,
	output wire [QUAN_SIZE-1:0] msg_out_6,
	output wire [QUAN_SIZE-1:0] msg_out_7,
	output wire [QUAN_SIZE-1:0] msg_out_8,
	output wire [QUAN_SIZE-1:0] msg_out_9,
	output wire [QUAN_SIZE-1:0] msg_out_10,
	output wire [QUAN_SIZE-1:0] msg_out_11,
	output wire [QUAN_SIZE-1:0] msg_out_12,
	output wire [QUAN_SIZE-1:0] msg_out_13,
	output wire [QUAN_SIZE-1:0] msg_out_14,
	output wire [QUAN_SIZE-1:0] msg_out_15,
	output wire [QUAN_SIZE-1:0] msg_out_16,
	output wire [QUAN_SIZE-1:0] msg_out_17,
	output wire [QUAN_SIZE-1:0] msg_out_18,
	output wire [QUAN_SIZE-1:0] msg_out_19,
	output wire [QUAN_SIZE-1:0] msg_out_20,
	output wire [QUAN_SIZE-1:0] msg_out_21,
	output wire [QUAN_SIZE-1:0] msg_out_22,
	output wire [QUAN_SIZE-1:0] msg_out_23,
	output wire [QUAN_SIZE-1:0] msg_out_24,
	output wire [QUAN_SIZE-1:0] msg_out_25,
	output wire [QUAN_SIZE-1:0] msg_out_26,
	output wire [QUAN_SIZE-1:0] msg_out_27,
	output wire [QUAN_SIZE-1:0] msg_out_28,
	output wire [QUAN_SIZE-1:0] msg_out_29,
	output wire [QUAN_SIZE-1:0] msg_out_30,
	output wire [QUAN_SIZE-1:0] msg_out_31,
	output wire [QUAN_SIZE-1:0] msg_out_32,
	output wire [QUAN_SIZE-1:0] msg_out_33,
	output wire [QUAN_SIZE-1:0] msg_out_34,
	output wire [QUAN_SIZE-1:0] msg_out_35,
	output wire [QUAN_SIZE-1:0] msg_out_36,
	output wire [QUAN_SIZE-1:0] msg_out_37,
	output wire [QUAN_SIZE-1:0] msg_out_38,
	output wire [QUAN_SIZE-1:0] msg_out_39,
	output wire [QUAN_SIZE-1:0] msg_out_40,
	output wire [QUAN_SIZE-1:0] msg_out_41,
	output wire [QUAN_SIZE-1:0] msg_out_42,
	output wire [QUAN_SIZE-1:0] msg_out_43,
	output wire [QUAN_SIZE-1:0] msg_out_44,
	output wire [QUAN_SIZE-1:0] msg_out_45,
	output wire [QUAN_SIZE-1:0] msg_out_46,
	output wire [QUAN_SIZE-1:0] msg_out_47,
	output wire [QUAN_SIZE-1:0] msg_out_48,
	output wire [QUAN_SIZE-1:0] msg_out_49,
	output wire [QUAN_SIZE-1:0] msg_out_50,
	output wire [QUAN_SIZE-1:0] msg_out_51,
	output wire [QUAN_SIZE-1:0] msg_out_52,
	output wire [QUAN_SIZE-1:0] msg_out_53,
	output wire [QUAN_SIZE-1:0] msg_out_54,
	output wire [QUAN_SIZE-1:0] msg_out_55,
	output wire [QUAN_SIZE-1:0] msg_out_56,
	output wire [QUAN_SIZE-1:0] msg_out_57,
	output wire [QUAN_SIZE-1:0] msg_out_58,
	output wire [QUAN_SIZE-1:0] msg_out_59,
	output wire [QUAN_SIZE-1:0] msg_out_60,
	output wire [QUAN_SIZE-1:0] msg_out_61,
	output wire [QUAN_SIZE-1:0] msg_out_62,
	output wire [QUAN_SIZE-1:0] msg_out_63,
	output wire [QUAN_SIZE-1:0] msg_out_64,
	output wire [QUAN_SIZE-1:0] msg_out_65,
	output wire [QUAN_SIZE-1:0] msg_out_66,
	output wire [QUAN_SIZE-1:0] msg_out_67,
	output wire [QUAN_SIZE-1:0] msg_out_68,
	output wire [QUAN_SIZE-1:0] msg_out_69,
	output wire [QUAN_SIZE-1:0] msg_out_70,
	output wire [QUAN_SIZE-1:0] msg_out_71,
	output wire [QUAN_SIZE-1:0] msg_out_72,
	output wire [QUAN_SIZE-1:0] msg_out_73,
	output wire [QUAN_SIZE-1:0] msg_out_74,
	output wire [QUAN_SIZE-1:0] msg_out_75,
	output wire [QUAN_SIZE-1:0] msg_out_76,
	output wire [QUAN_SIZE-1:0] msg_out_77,
	output wire [QUAN_SIZE-1:0] msg_out_78,
	output wire [QUAN_SIZE-1:0] msg_out_79,
	output wire [QUAN_SIZE-1:0] msg_out_80,
	output wire [QUAN_SIZE-1:0] msg_out_81,
	output wire [QUAN_SIZE-1:0] msg_out_82,
	output wire [QUAN_SIZE-1:0] msg_out_83,
	output wire [QUAN_SIZE-1:0] msg_out_84,
	output wire [QUAN_SIZE-1:0] msg_out_85,
	output wire [QUAN_SIZE-1:0] msg_out_86,
	output wire [QUAN_SIZE-1:0] msg_out_87,
	output wire [QUAN_SIZE-1:0] msg_out_88,
	output wire [QUAN_SIZE-1:0] msg_out_89,
	output wire [QUAN_SIZE-1:0] msg_out_90,
	output wire [QUAN_SIZE-1:0] msg_out_91,
	output wire [QUAN_SIZE-1:0] msg_out_92,
	output wire [QUAN_SIZE-1:0] msg_out_93,
	output wire [QUAN_SIZE-1:0] msg_out_94,
	output wire [QUAN_SIZE-1:0] msg_out_95,
	output wire [QUAN_SIZE-1:0] msg_out_96,
	output wire [QUAN_SIZE-1:0] msg_out_97,
	output wire [QUAN_SIZE-1:0] msg_out_98,
	output wire [QUAN_SIZE-1:0] msg_out_99,
	output wire [QUAN_SIZE-1:0] msg_out_100,
	output wire [QUAN_SIZE-1:0] msg_out_101,
	output wire [QUAN_SIZE-1:0] msg_out_102,
	output wire [QUAN_SIZE-1:0] msg_out_103,
	output wire [QUAN_SIZE-1:0] msg_out_104,
	output wire [QUAN_SIZE-1:0] msg_out_105,
	output wire [QUAN_SIZE-1:0] msg_out_106,
	output wire [QUAN_SIZE-1:0] msg_out_107,
	output wire [QUAN_SIZE-1:0] msg_out_108,
	output wire [QUAN_SIZE-1:0] msg_out_109,
	output wire [QUAN_SIZE-1:0] msg_out_110,
	output wire [QUAN_SIZE-1:0] msg_out_111,
	output wire [QUAN_SIZE-1:0] msg_out_112,
	output wire [QUAN_SIZE-1:0] msg_out_113,
	output wire [QUAN_SIZE-1:0] msg_out_114,
	output wire [QUAN_SIZE-1:0] msg_out_115,
	output wire [QUAN_SIZE-1:0] msg_out_116,
	output wire [QUAN_SIZE-1:0] msg_out_117,
	output wire [QUAN_SIZE-1:0] msg_out_118,
	output wire [QUAN_SIZE-1:0] msg_out_119,
	output wire [QUAN_SIZE-1:0] msg_out_120,
	output wire [QUAN_SIZE-1:0] msg_out_121,
	output wire [QUAN_SIZE-1:0] msg_out_122,
	output wire [QUAN_SIZE-1:0] msg_out_123,
	output wire [QUAN_SIZE-1:0] msg_out_124,
	output wire [QUAN_SIZE-1:0] msg_out_125,
	output wire [QUAN_SIZE-1:0] msg_out_126,
	output wire [QUAN_SIZE-1:0] msg_out_127,
	output wire [QUAN_SIZE-1:0] msg_out_128,
	output wire [QUAN_SIZE-1:0] msg_out_129,
	output wire [QUAN_SIZE-1:0] msg_out_130,
	output wire [QUAN_SIZE-1:0] msg_out_131,
	output wire [QUAN_SIZE-1:0] msg_out_132,
	output wire [QUAN_SIZE-1:0] msg_out_133,
	output wire [QUAN_SIZE-1:0] msg_out_134,
	output wire [QUAN_SIZE-1:0] msg_out_135,
	output wire [QUAN_SIZE-1:0] msg_out_136,
	output wire [QUAN_SIZE-1:0] msg_out_137,
	output wire [QUAN_SIZE-1:0] msg_out_138,
	output wire [QUAN_SIZE-1:0] msg_out_139,
	output wire [QUAN_SIZE-1:0] msg_out_140,
	output wire [QUAN_SIZE-1:0] msg_out_141,
	output wire [QUAN_SIZE-1:0] msg_out_142,
	output wire [QUAN_SIZE-1:0] msg_out_143,
	output wire [QUAN_SIZE-1:0] msg_out_144,
	output wire [QUAN_SIZE-1:0] msg_out_145,
	output wire [QUAN_SIZE-1:0] msg_out_146,
	output wire [QUAN_SIZE-1:0] msg_out_147,
	output wire [QUAN_SIZE-1:0] msg_out_148,
	output wire [QUAN_SIZE-1:0] msg_out_149,
	output wire [QUAN_SIZE-1:0] msg_out_150,
	output wire [QUAN_SIZE-1:0] msg_out_151,
	output wire [QUAN_SIZE-1:0] msg_out_152,
	output wire [QUAN_SIZE-1:0] msg_out_153,
	output wire [QUAN_SIZE-1:0] msg_out_154,
	output wire [QUAN_SIZE-1:0] msg_out_155,
	output wire [QUAN_SIZE-1:0] msg_out_156,
	output wire [QUAN_SIZE-1:0] msg_out_157,
	output wire [QUAN_SIZE-1:0] msg_out_158,
	output wire [QUAN_SIZE-1:0] msg_out_159,
	output wire [QUAN_SIZE-1:0] msg_out_160,
	output wire [QUAN_SIZE-1:0] msg_out_161,
	output wire [QUAN_SIZE-1:0] msg_out_162,
	output wire [QUAN_SIZE-1:0] msg_out_163,
	output wire [QUAN_SIZE-1:0] msg_out_164,
	output wire [QUAN_SIZE-1:0] msg_out_165,
	output wire [QUAN_SIZE-1:0] msg_out_166,
	output wire [QUAN_SIZE-1:0] msg_out_167,
	output wire [QUAN_SIZE-1:0] msg_out_168,
	output wire [QUAN_SIZE-1:0] msg_out_169,
	output wire [QUAN_SIZE-1:0] msg_out_170,
	output wire [QUAN_SIZE-1:0] msg_out_171,
	output wire [QUAN_SIZE-1:0] msg_out_172,
	output wire [QUAN_SIZE-1:0] msg_out_173,
	output wire [QUAN_SIZE-1:0] msg_out_174,
	output wire [QUAN_SIZE-1:0] msg_out_175,
	output wire [QUAN_SIZE-1:0] msg_out_176,
	output wire [QUAN_SIZE-1:0] msg_out_177,
	output wire [QUAN_SIZE-1:0] msg_out_178,
	output wire [QUAN_SIZE-1:0] msg_out_179,
	output wire [QUAN_SIZE-1:0] msg_out_180,
	output wire [QUAN_SIZE-1:0] msg_out_181,
	output wire [QUAN_SIZE-1:0] msg_out_182,
	output wire [QUAN_SIZE-1:0] msg_out_183,
	output wire [QUAN_SIZE-1:0] msg_out_184,
	output wire [QUAN_SIZE-1:0] msg_out_185,
	output wire [QUAN_SIZE-1:0] msg_out_186,
	output wire [QUAN_SIZE-1:0] msg_out_187,
	output wire [QUAN_SIZE-1:0] msg_out_188,
	output wire [QUAN_SIZE-1:0] msg_out_189,
	output wire [QUAN_SIZE-1:0] msg_out_190,
	output wire [QUAN_SIZE-1:0] msg_out_191,
	output wire [QUAN_SIZE-1:0] msg_out_192,
	output wire [QUAN_SIZE-1:0] msg_out_193,
	output wire [QUAN_SIZE-1:0] msg_out_194,
	output wire [QUAN_SIZE-1:0] msg_out_195,
	output wire [QUAN_SIZE-1:0] msg_out_196,
	output wire [QUAN_SIZE-1:0] msg_out_197,
	output wire [QUAN_SIZE-1:0] msg_out_198,
	output wire [QUAN_SIZE-1:0] msg_out_199,
	output wire [QUAN_SIZE-1:0] msg_out_200,
	output wire [QUAN_SIZE-1:0] msg_out_201,
	output wire [QUAN_SIZE-1:0] msg_out_202,
	output wire [QUAN_SIZE-1:0] msg_out_203,
	output wire [QUAN_SIZE-1:0] msg_out_204,
	output wire [QUAN_SIZE-1:0] msg_out_205,
	output wire [QUAN_SIZE-1:0] msg_out_206,
	output wire [QUAN_SIZE-1:0] msg_out_207,
	output wire [QUAN_SIZE-1:0] msg_out_208,
	output wire [QUAN_SIZE-1:0] msg_out_209,
	output wire [QUAN_SIZE-1:0] msg_out_210,
	output wire [QUAN_SIZE-1:0] msg_out_211,
	output wire [QUAN_SIZE-1:0] msg_out_212,
	output wire [QUAN_SIZE-1:0] msg_out_213,
	output wire [QUAN_SIZE-1:0] msg_out_214,
	output wire [QUAN_SIZE-1:0] msg_out_215,
	output wire [QUAN_SIZE-1:0] msg_out_216,
	output wire [QUAN_SIZE-1:0] msg_out_217,
	output wire [QUAN_SIZE-1:0] msg_out_218,
	output wire [QUAN_SIZE-1:0] msg_out_219,
	output wire [QUAN_SIZE-1:0] msg_out_220,
	output wire [QUAN_SIZE-1:0] msg_out_221,
	output wire [QUAN_SIZE-1:0] msg_out_222,
	output wire [QUAN_SIZE-1:0] msg_out_223,
	output wire [QUAN_SIZE-1:0] msg_out_224,
	output wire [QUAN_SIZE-1:0] msg_out_225,
	output wire [QUAN_SIZE-1:0] msg_out_226,
	output wire [QUAN_SIZE-1:0] msg_out_227,
	output wire [QUAN_SIZE-1:0] msg_out_228,
	output wire [QUAN_SIZE-1:0] msg_out_229,
	output wire [QUAN_SIZE-1:0] msg_out_230,
	output wire [QUAN_SIZE-1:0] msg_out_231,
	output wire [QUAN_SIZE-1:0] msg_out_232,
	output wire [QUAN_SIZE-1:0] msg_out_233,
	output wire [QUAN_SIZE-1:0] msg_out_234,
	output wire [QUAN_SIZE-1:0] msg_out_235,
	output wire [QUAN_SIZE-1:0] msg_out_236,
	output wire [QUAN_SIZE-1:0] msg_out_237,
	output wire [QUAN_SIZE-1:0] msg_out_238,
	output wire [QUAN_SIZE-1:0] msg_out_239,
	output wire [QUAN_SIZE-1:0] msg_out_240,
	output wire [QUAN_SIZE-1:0] msg_out_241,
	output wire [QUAN_SIZE-1:0] msg_out_242,
	output wire [QUAN_SIZE-1:0] msg_out_243,
	output wire [QUAN_SIZE-1:0] msg_out_244,
	output wire [QUAN_SIZE-1:0] msg_out_245,
	output wire [QUAN_SIZE-1:0] msg_out_246,
	output wire [QUAN_SIZE-1:0] msg_out_247,
	output wire [QUAN_SIZE-1:0] msg_out_248,
	output wire [QUAN_SIZE-1:0] msg_out_249,
	output wire [QUAN_SIZE-1:0] msg_out_250,
	output wire [QUAN_SIZE-1:0] msg_out_251,
	output wire [QUAN_SIZE-1:0] msg_out_252,
	output wire [QUAN_SIZE-1:0] msg_out_253,
	output wire [QUAN_SIZE-1:0] msg_out_254,

	input wire [QUAN_SIZE-1:0] msg_in_0,
	input wire [QUAN_SIZE-1:0] msg_in_1,
	input wire [QUAN_SIZE-1:0] msg_in_2,
	input wire [QUAN_SIZE-1:0] msg_in_3,
	input wire [QUAN_SIZE-1:0] msg_in_4,
	input wire [QUAN_SIZE-1:0] msg_in_5,
	input wire [QUAN_SIZE-1:0] msg_in_6,
	input wire [QUAN_SIZE-1:0] msg_in_7,
	input wire [QUAN_SIZE-1:0] msg_in_8,
	input wire [QUAN_SIZE-1:0] msg_in_9,
	input wire [QUAN_SIZE-1:0] msg_in_10,
	input wire [QUAN_SIZE-1:0] msg_in_11,
	input wire [QUAN_SIZE-1:0] msg_in_12,
	input wire [QUAN_SIZE-1:0] msg_in_13,
	input wire [QUAN_SIZE-1:0] msg_in_14,
	input wire [QUAN_SIZE-1:0] msg_in_15,
	input wire [QUAN_SIZE-1:0] msg_in_16,
	input wire [QUAN_SIZE-1:0] msg_in_17,
	input wire [QUAN_SIZE-1:0] msg_in_18,
	input wire [QUAN_SIZE-1:0] msg_in_19,
	input wire [QUAN_SIZE-1:0] msg_in_20,
	input wire [QUAN_SIZE-1:0] msg_in_21,
	input wire [QUAN_SIZE-1:0] msg_in_22,
	input wire [QUAN_SIZE-1:0] msg_in_23,
	input wire [QUAN_SIZE-1:0] msg_in_24,
	input wire [QUAN_SIZE-1:0] msg_in_25,
	input wire [QUAN_SIZE-1:0] msg_in_26,
	input wire [QUAN_SIZE-1:0] msg_in_27,
	input wire [QUAN_SIZE-1:0] msg_in_28,
	input wire [QUAN_SIZE-1:0] msg_in_29,
	input wire [QUAN_SIZE-1:0] msg_in_30,
	input wire [QUAN_SIZE-1:0] msg_in_31,
	input wire [QUAN_SIZE-1:0] msg_in_32,
	input wire [QUAN_SIZE-1:0] msg_in_33,
	input wire [QUAN_SIZE-1:0] msg_in_34,
	input wire [QUAN_SIZE-1:0] msg_in_35,
	input wire [QUAN_SIZE-1:0] msg_in_36,
	input wire [QUAN_SIZE-1:0] msg_in_37,
	input wire [QUAN_SIZE-1:0] msg_in_38,
	input wire [QUAN_SIZE-1:0] msg_in_39,
	input wire [QUAN_SIZE-1:0] msg_in_40,
	input wire [QUAN_SIZE-1:0] msg_in_41,
	input wire [QUAN_SIZE-1:0] msg_in_42,
	input wire [QUAN_SIZE-1:0] msg_in_43,
	input wire [QUAN_SIZE-1:0] msg_in_44,
	input wire [QUAN_SIZE-1:0] msg_in_45,
	input wire [QUAN_SIZE-1:0] msg_in_46,
	input wire [QUAN_SIZE-1:0] msg_in_47,
	input wire [QUAN_SIZE-1:0] msg_in_48,
	input wire [QUAN_SIZE-1:0] msg_in_49,
	input wire [QUAN_SIZE-1:0] msg_in_50,
	input wire [QUAN_SIZE-1:0] msg_in_51,
	input wire [QUAN_SIZE-1:0] msg_in_52,
	input wire [QUAN_SIZE-1:0] msg_in_53,
	input wire [QUAN_SIZE-1:0] msg_in_54,
	input wire [QUAN_SIZE-1:0] msg_in_55,
	input wire [QUAN_SIZE-1:0] msg_in_56,
	input wire [QUAN_SIZE-1:0] msg_in_57,
	input wire [QUAN_SIZE-1:0] msg_in_58,
	input wire [QUAN_SIZE-1:0] msg_in_59,
	input wire [QUAN_SIZE-1:0] msg_in_60,
	input wire [QUAN_SIZE-1:0] msg_in_61,
	input wire [QUAN_SIZE-1:0] msg_in_62,
	input wire [QUAN_SIZE-1:0] msg_in_63,
	input wire [QUAN_SIZE-1:0] msg_in_64,
	input wire [QUAN_SIZE-1:0] msg_in_65,
	input wire [QUAN_SIZE-1:0] msg_in_66,
	input wire [QUAN_SIZE-1:0] msg_in_67,
	input wire [QUAN_SIZE-1:0] msg_in_68,
	input wire [QUAN_SIZE-1:0] msg_in_69,
	input wire [QUAN_SIZE-1:0] msg_in_70,
	input wire [QUAN_SIZE-1:0] msg_in_71,
	input wire [QUAN_SIZE-1:0] msg_in_72,
	input wire [QUAN_SIZE-1:0] msg_in_73,
	input wire [QUAN_SIZE-1:0] msg_in_74,
	input wire [QUAN_SIZE-1:0] msg_in_75,
	input wire [QUAN_SIZE-1:0] msg_in_76,
	input wire [QUAN_SIZE-1:0] msg_in_77,
	input wire [QUAN_SIZE-1:0] msg_in_78,
	input wire [QUAN_SIZE-1:0] msg_in_79,
	input wire [QUAN_SIZE-1:0] msg_in_80,
	input wire [QUAN_SIZE-1:0] msg_in_81,
	input wire [QUAN_SIZE-1:0] msg_in_82,
	input wire [QUAN_SIZE-1:0] msg_in_83,
	input wire [QUAN_SIZE-1:0] msg_in_84,
	input wire [QUAN_SIZE-1:0] msg_in_85,
	input wire [QUAN_SIZE-1:0] msg_in_86,
	input wire [QUAN_SIZE-1:0] msg_in_87,
	input wire [QUAN_SIZE-1:0] msg_in_88,
	input wire [QUAN_SIZE-1:0] msg_in_89,
	input wire [QUAN_SIZE-1:0] msg_in_90,
	input wire [QUAN_SIZE-1:0] msg_in_91,
	input wire [QUAN_SIZE-1:0] msg_in_92,
	input wire [QUAN_SIZE-1:0] msg_in_93,
	input wire [QUAN_SIZE-1:0] msg_in_94,
	input wire [QUAN_SIZE-1:0] msg_in_95,
	input wire [QUAN_SIZE-1:0] msg_in_96,
	input wire [QUAN_SIZE-1:0] msg_in_97,
	input wire [QUAN_SIZE-1:0] msg_in_98,
	input wire [QUAN_SIZE-1:0] msg_in_99,
	input wire [QUAN_SIZE-1:0] msg_in_100,
	input wire [QUAN_SIZE-1:0] msg_in_101,
	input wire [QUAN_SIZE-1:0] msg_in_102,
	input wire [QUAN_SIZE-1:0] msg_in_103,
	input wire [QUAN_SIZE-1:0] msg_in_104,
	input wire [QUAN_SIZE-1:0] msg_in_105,
	input wire [QUAN_SIZE-1:0] msg_in_106,
	input wire [QUAN_SIZE-1:0] msg_in_107,
	input wire [QUAN_SIZE-1:0] msg_in_108,
	input wire [QUAN_SIZE-1:0] msg_in_109,
	input wire [QUAN_SIZE-1:0] msg_in_110,
	input wire [QUAN_SIZE-1:0] msg_in_111,
	input wire [QUAN_SIZE-1:0] msg_in_112,
	input wire [QUAN_SIZE-1:0] msg_in_113,
	input wire [QUAN_SIZE-1:0] msg_in_114,
	input wire [QUAN_SIZE-1:0] msg_in_115,
	input wire [QUAN_SIZE-1:0] msg_in_116,
	input wire [QUAN_SIZE-1:0] msg_in_117,
	input wire [QUAN_SIZE-1:0] msg_in_118,
	input wire [QUAN_SIZE-1:0] msg_in_119,
	input wire [QUAN_SIZE-1:0] msg_in_120,
	input wire [QUAN_SIZE-1:0] msg_in_121,
	input wire [QUAN_SIZE-1:0] msg_in_122,
	input wire [QUAN_SIZE-1:0] msg_in_123,
	input wire [QUAN_SIZE-1:0] msg_in_124,
	input wire [QUAN_SIZE-1:0] msg_in_125,
	input wire [QUAN_SIZE-1:0] msg_in_126,
	input wire [QUAN_SIZE-1:0] msg_in_127,
	input wire [QUAN_SIZE-1:0] msg_in_128,
	input wire [QUAN_SIZE-1:0] msg_in_129,
	input wire [QUAN_SIZE-1:0] msg_in_130,
	input wire [QUAN_SIZE-1:0] msg_in_131,
	input wire [QUAN_SIZE-1:0] msg_in_132,
	input wire [QUAN_SIZE-1:0] msg_in_133,
	input wire [QUAN_SIZE-1:0] msg_in_134,
	input wire [QUAN_SIZE-1:0] msg_in_135,
	input wire [QUAN_SIZE-1:0] msg_in_136,
	input wire [QUAN_SIZE-1:0] msg_in_137,
	input wire [QUAN_SIZE-1:0] msg_in_138,
	input wire [QUAN_SIZE-1:0] msg_in_139,
	input wire [QUAN_SIZE-1:0] msg_in_140,
	input wire [QUAN_SIZE-1:0] msg_in_141,
	input wire [QUAN_SIZE-1:0] msg_in_142,
	input wire [QUAN_SIZE-1:0] msg_in_143,
	input wire [QUAN_SIZE-1:0] msg_in_144,
	input wire [QUAN_SIZE-1:0] msg_in_145,
	input wire [QUAN_SIZE-1:0] msg_in_146,
	input wire [QUAN_SIZE-1:0] msg_in_147,
	input wire [QUAN_SIZE-1:0] msg_in_148,
	input wire [QUAN_SIZE-1:0] msg_in_149,
	input wire [QUAN_SIZE-1:0] msg_in_150,
	input wire [QUAN_SIZE-1:0] msg_in_151,
	input wire [QUAN_SIZE-1:0] msg_in_152,
	input wire [QUAN_SIZE-1:0] msg_in_153,
	input wire [QUAN_SIZE-1:0] msg_in_154,
	input wire [QUAN_SIZE-1:0] msg_in_155,
	input wire [QUAN_SIZE-1:0] msg_in_156,
	input wire [QUAN_SIZE-1:0] msg_in_157,
	input wire [QUAN_SIZE-1:0] msg_in_158,
	input wire [QUAN_SIZE-1:0] msg_in_159,
	input wire [QUAN_SIZE-1:0] msg_in_160,
	input wire [QUAN_SIZE-1:0] msg_in_161,
	input wire [QUAN_SIZE-1:0] msg_in_162,
	input wire [QUAN_SIZE-1:0] msg_in_163,
	input wire [QUAN_SIZE-1:0] msg_in_164,
	input wire [QUAN_SIZE-1:0] msg_in_165,
	input wire [QUAN_SIZE-1:0] msg_in_166,
	input wire [QUAN_SIZE-1:0] msg_in_167,
	input wire [QUAN_SIZE-1:0] msg_in_168,
	input wire [QUAN_SIZE-1:0] msg_in_169,
	input wire [QUAN_SIZE-1:0] msg_in_170,
	input wire [QUAN_SIZE-1:0] msg_in_171,
	input wire [QUAN_SIZE-1:0] msg_in_172,
	input wire [QUAN_SIZE-1:0] msg_in_173,
	input wire [QUAN_SIZE-1:0] msg_in_174,
	input wire [QUAN_SIZE-1:0] msg_in_175,
	input wire [QUAN_SIZE-1:0] msg_in_176,
	input wire [QUAN_SIZE-1:0] msg_in_177,
	input wire [QUAN_SIZE-1:0] msg_in_178,
	input wire [QUAN_SIZE-1:0] msg_in_179,
	input wire [QUAN_SIZE-1:0] msg_in_180,
	input wire [QUAN_SIZE-1:0] msg_in_181,
	input wire [QUAN_SIZE-1:0] msg_in_182,
	input wire [QUAN_SIZE-1:0] msg_in_183,
	input wire [QUAN_SIZE-1:0] msg_in_184,
	input wire [QUAN_SIZE-1:0] msg_in_185,
	input wire [QUAN_SIZE-1:0] msg_in_186,
	input wire [QUAN_SIZE-1:0] msg_in_187,
	input wire [QUAN_SIZE-1:0] msg_in_188,
	input wire [QUAN_SIZE-1:0] msg_in_189,
	input wire [QUAN_SIZE-1:0] msg_in_190,
	input wire [QUAN_SIZE-1:0] msg_in_191,
	input wire [QUAN_SIZE-1:0] msg_in_192,
	input wire [QUAN_SIZE-1:0] msg_in_193,
	input wire [QUAN_SIZE-1:0] msg_in_194,
	input wire [QUAN_SIZE-1:0] msg_in_195,
	input wire [QUAN_SIZE-1:0] msg_in_196,
	input wire [QUAN_SIZE-1:0] msg_in_197,
	input wire [QUAN_SIZE-1:0] msg_in_198,
	input wire [QUAN_SIZE-1:0] msg_in_199,
	input wire [QUAN_SIZE-1:0] msg_in_200,
	input wire [QUAN_SIZE-1:0] msg_in_201,
	input wire [QUAN_SIZE-1:0] msg_in_202,
	input wire [QUAN_SIZE-1:0] msg_in_203,
	input wire [QUAN_SIZE-1:0] msg_in_204,
	input wire [QUAN_SIZE-1:0] msg_in_205,
	input wire [QUAN_SIZE-1:0] msg_in_206,
	input wire [QUAN_SIZE-1:0] msg_in_207,
	input wire [QUAN_SIZE-1:0] msg_in_208,
	input wire [QUAN_SIZE-1:0] msg_in_209,
	input wire [QUAN_SIZE-1:0] msg_in_210,
	input wire [QUAN_SIZE-1:0] msg_in_211,
	input wire [QUAN_SIZE-1:0] msg_in_212,
	input wire [QUAN_SIZE-1:0] msg_in_213,
	input wire [QUAN_SIZE-1:0] msg_in_214,
	input wire [QUAN_SIZE-1:0] msg_in_215,
	input wire [QUAN_SIZE-1:0] msg_in_216,
	input wire [QUAN_SIZE-1:0] msg_in_217,
	input wire [QUAN_SIZE-1:0] msg_in_218,
	input wire [QUAN_SIZE-1:0] msg_in_219,
	input wire [QUAN_SIZE-1:0] msg_in_220,
	input wire [QUAN_SIZE-1:0] msg_in_221,
	input wire [QUAN_SIZE-1:0] msg_in_222,
	input wire [QUAN_SIZE-1:0] msg_in_223,
	input wire [QUAN_SIZE-1:0] msg_in_224,
	input wire [QUAN_SIZE-1:0] msg_in_225,
	input wire [QUAN_SIZE-1:0] msg_in_226,
	input wire [QUAN_SIZE-1:0] msg_in_227,
	input wire [QUAN_SIZE-1:0] msg_in_228,
	input wire [QUAN_SIZE-1:0] msg_in_229,
	input wire [QUAN_SIZE-1:0] msg_in_230,
	input wire [QUAN_SIZE-1:0] msg_in_231,
	input wire [QUAN_SIZE-1:0] msg_in_232,
	input wire [QUAN_SIZE-1:0] msg_in_233,
	input wire [QUAN_SIZE-1:0] msg_in_234,
	input wire [QUAN_SIZE-1:0] msg_in_235,
	input wire [QUAN_SIZE-1:0] msg_in_236,
	input wire [QUAN_SIZE-1:0] msg_in_237,
	input wire [QUAN_SIZE-1:0] msg_in_238,
	input wire [QUAN_SIZE-1:0] msg_in_239,
	input wire [QUAN_SIZE-1:0] msg_in_240,
	input wire [QUAN_SIZE-1:0] msg_in_241,
	input wire [QUAN_SIZE-1:0] msg_in_242,
	input wire [QUAN_SIZE-1:0] msg_in_243,
	input wire [QUAN_SIZE-1:0] msg_in_244,
	input wire [QUAN_SIZE-1:0] msg_in_245,
	input wire [QUAN_SIZE-1:0] msg_in_246,
	input wire [QUAN_SIZE-1:0] msg_in_247,
	input wire [QUAN_SIZE-1:0] msg_in_248,
	input wire [QUAN_SIZE-1:0] msg_in_249,
	input wire [QUAN_SIZE-1:0] msg_in_250,
	input wire [QUAN_SIZE-1:0] msg_in_251,
	input wire [QUAN_SIZE-1:0] msg_in_252,
	input wire [QUAN_SIZE-1:0] msg_in_253,
	input wire [QUAN_SIZE-1:0] msg_in_254,

	input wire [LAYER_NUM-1:0] layer_status,
	input wire first_row_chunk,
	input wire sys_clk,
	input wire rstn
);

/////////////////////////////////////////////////////////////////////////////////////////////
// Main structure of Page Alignment Mechanism
wire [1:0] sub_4_circular_delay_cmd_1_4;
assign sub_4_circular_delay_cmd_1_4 = ((layer_status[0] == 1'b1 || layer_status[2] == 1'b1) && first_row_chunk == 1'b1) ? 2'b10 : (layer_status[1] == 1'b1) ? 2'b01 : 2'b00;
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u77 (.align_out (msg_out_77), .align_target_in (msg_in_77), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u78 (.align_out (msg_out_78), .align_target_in (msg_in_78), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u79 (.align_out (msg_out_79), .align_target_in (msg_in_79), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u80 (.align_out (msg_out_80), .align_target_in (msg_in_80), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u81 (.align_out (msg_out_81), .align_target_in (msg_in_81), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u82 (.align_out (msg_out_82), .align_target_in (msg_in_82), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u83 (.align_out (msg_out_83), .align_target_in (msg_in_83), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u84 (.align_out (msg_out_84), .align_target_in (msg_in_84), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u85 (.align_out (msg_out_85), .align_target_in (msg_in_85), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u86 (.align_out (msg_out_86), .align_target_in (msg_in_86), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u87 (.align_out (msg_out_87), .align_target_in (msg_in_87), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u88 (.align_out (msg_out_88), .align_target_in (msg_in_88), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u89 (.align_out (msg_out_89), .align_target_in (msg_in_89), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u90 (.align_out (msg_out_90), .align_target_in (msg_in_90), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u91 (.align_out (msg_out_91), .align_target_in (msg_in_91), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u92 (.align_out (msg_out_92), .align_target_in (msg_in_92), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u93 (.align_out (msg_out_93), .align_target_in (msg_in_93), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u94 (.align_out (msg_out_94), .align_target_in (msg_in_94), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u95 (.align_out (msg_out_95), .align_target_in (msg_in_95), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u96 (.align_out (msg_out_96), .align_target_in (msg_in_96), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u97 (.align_out (msg_out_97), .align_target_in (msg_in_97), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u98 (.align_out (msg_out_98), .align_target_in (msg_in_98), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u99 (.align_out (msg_out_99), .align_target_in (msg_in_99), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u100 (.align_out (msg_out_100), .align_target_in (msg_in_100), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u101 (.align_out (msg_out_101), .align_target_in (msg_in_101), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u102 (.align_out (msg_out_102), .align_target_in (msg_in_102), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u103 (.align_out (msg_out_103), .align_target_in (msg_in_103), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u104 (.align_out (msg_out_104), .align_target_in (msg_in_104), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u105 (.align_out (msg_out_105), .align_target_in (msg_in_105), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u106 (.align_out (msg_out_106), .align_target_in (msg_in_106), .delay_cmd(sub_4_circular_delay_cmd_1_4), .sys_clk(sys_clk), .rstn(rstn));
wire [1:0] sub_4_circular_delay_cmd_5_0;
assign sub_4_circular_delay_cmd_5_0 = (layer_status[0] == 1'b1 && first_row_chunk == 1'b1) ? 2'b10 : (layer_status[1] == 1'b1 || layer_status[2] == 1'b1) ? 2'b01 : 2'b00;
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u71 (.align_out (msg_out_71), .align_target_in (msg_in_71), .delay_cmd(sub_4_circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u72 (.align_out (msg_out_72), .align_target_in (msg_in_72), .delay_cmd(sub_4_circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u73 (.align_out (msg_out_73), .align_target_in (msg_in_73), .delay_cmd(sub_4_circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u74 (.align_out (msg_out_74), .align_target_in (msg_in_74), .delay_cmd(sub_4_circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u75 (.align_out (msg_out_75), .align_target_in (msg_in_75), .delay_cmd(sub_4_circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u76 (.align_out (msg_out_76), .align_target_in (msg_in_76), .delay_cmd(sub_4_circular_delay_cmd_5_0), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u0(.align_out(msg_out_0), .align_target_in (msg_in_0), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u1(.align_out(msg_out_1), .align_target_in (msg_in_1), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u2(.align_out(msg_out_2), .align_target_in (msg_in_2), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u3(.align_out(msg_out_3), .align_target_in (msg_in_3), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u4(.align_out(msg_out_4), .align_target_in (msg_in_4), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u5(.align_out(msg_out_5), .align_target_in (msg_in_5), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u6(.align_out(msg_out_6), .align_target_in (msg_in_6), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u7(.align_out(msg_out_7), .align_target_in (msg_in_7), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u8(.align_out(msg_out_8), .align_target_in (msg_in_8), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u9(.align_out(msg_out_9), .align_target_in (msg_in_9), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u10(.align_out(msg_out_10), .align_target_in (msg_in_10), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u11(.align_out(msg_out_11), .align_target_in (msg_in_11), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u12(.align_out(msg_out_12), .align_target_in (msg_in_12), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u13(.align_out(msg_out_13), .align_target_in (msg_in_13), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u14(.align_out(msg_out_14), .align_target_in (msg_in_14), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u15(.align_out(msg_out_15), .align_target_in (msg_in_15), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u16(.align_out(msg_out_16), .align_target_in (msg_in_16), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u17(.align_out(msg_out_17), .align_target_in (msg_in_17), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u18(.align_out(msg_out_18), .align_target_in (msg_in_18), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u19(.align_out(msg_out_19), .align_target_in (msg_in_19), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u20(.align_out(msg_out_20), .align_target_in (msg_in_20), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u21(.align_out(msg_out_21), .align_target_in (msg_in_21), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u22(.align_out(msg_out_22), .align_target_in (msg_in_22), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u23(.align_out(msg_out_23), .align_target_in (msg_in_23), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u24(.align_out(msg_out_24), .align_target_in (msg_in_24), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u25(.align_out(msg_out_25), .align_target_in (msg_in_25), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u26(.align_out(msg_out_26), .align_target_in (msg_in_26), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u27(.align_out(msg_out_27), .align_target_in (msg_in_27), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u28(.align_out(msg_out_28), .align_target_in (msg_in_28), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u29(.align_out(msg_out_29), .align_target_in (msg_in_29), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u30(.align_out(msg_out_30), .align_target_in (msg_in_30), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u31(.align_out(msg_out_31), .align_target_in (msg_in_31), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u32(.align_out(msg_out_32), .align_target_in (msg_in_32), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u33(.align_out(msg_out_33), .align_target_in (msg_in_33), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u34(.align_out(msg_out_34), .align_target_in (msg_in_34), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u35(.align_out(msg_out_35), .align_target_in (msg_in_35), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u36(.align_out(msg_out_36), .align_target_in (msg_in_36), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u37(.align_out(msg_out_37), .align_target_in (msg_in_37), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u38(.align_out(msg_out_38), .align_target_in (msg_in_38), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u39(.align_out(msg_out_39), .align_target_in (msg_in_39), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u40(.align_out(msg_out_40), .align_target_in (msg_in_40), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u41(.align_out(msg_out_41), .align_target_in (msg_in_41), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u42(.align_out(msg_out_42), .align_target_in (msg_in_42), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u43(.align_out(msg_out_43), .align_target_in (msg_in_43), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u44(.align_out(msg_out_44), .align_target_in (msg_in_44), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u45(.align_out(msg_out_45), .align_target_in (msg_in_45), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u46(.align_out(msg_out_46), .align_target_in (msg_in_46), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u47(.align_out(msg_out_47), .align_target_in (msg_in_47), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u48(.align_out(msg_out_48), .align_target_in (msg_in_48), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u49(.align_out(msg_out_49), .align_target_in (msg_in_49), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u50(.align_out(msg_out_50), .align_target_in (msg_in_50), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u51(.align_out(msg_out_51), .align_target_in (msg_in_51), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u52(.align_out(msg_out_52), .align_target_in (msg_in_52), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u53(.align_out(msg_out_53), .align_target_in (msg_in_53), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u54(.align_out(msg_out_54), .align_target_in (msg_in_54), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u55(.align_out(msg_out_55), .align_target_in (msg_in_55), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u56(.align_out(msg_out_56), .align_target_in (msg_in_56), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u57(.align_out(msg_out_57), .align_target_in (msg_in_57), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u58(.align_out(msg_out_58), .align_target_in (msg_in_58), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u59(.align_out(msg_out_59), .align_target_in (msg_in_59), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u60(.align_out(msg_out_60), .align_target_in (msg_in_60), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u61(.align_out(msg_out_61), .align_target_in (msg_in_61), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u62(.align_out(msg_out_62), .align_target_in (msg_in_62), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u63(.align_out(msg_out_63), .align_target_in (msg_in_63), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u64(.align_out(msg_out_64), .align_target_in (msg_in_64), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u65(.align_out(msg_out_65), .align_target_in (msg_in_65), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u66(.align_out(msg_out_66), .align_target_in (msg_in_66), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u67(.align_out(msg_out_67), .align_target_in (msg_in_67), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u68(.align_out(msg_out_68), .align_target_in (msg_in_68), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u69(.align_out(msg_out_69), .align_target_in (msg_in_69), .sys_clk(sys_clk), .rstn(rstn));
page_align_depth_2 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u70(.align_out(msg_out_70), .align_target_in (msg_in_70), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u107 (.align_out (msg_out_107), .align_target_in (msg_in_107), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u108 (.align_out (msg_out_108), .align_target_in (msg_in_108), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u109 (.align_out (msg_out_109), .align_target_in (msg_in_109), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u110 (.align_out (msg_out_110), .align_target_in (msg_in_110), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u111 (.align_out (msg_out_111), .align_target_in (msg_in_111), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u112 (.align_out (msg_out_112), .align_target_in (msg_in_112), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u113 (.align_out (msg_out_113), .align_target_in (msg_in_113), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u114 (.align_out (msg_out_114), .align_target_in (msg_in_114), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u115 (.align_out (msg_out_115), .align_target_in (msg_in_115), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u116 (.align_out (msg_out_116), .align_target_in (msg_in_116), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u117 (.align_out (msg_out_117), .align_target_in (msg_in_117), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u118 (.align_out (msg_out_118), .align_target_in (msg_in_118), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u119 (.align_out (msg_out_119), .align_target_in (msg_in_119), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u120 (.align_out (msg_out_120), .align_target_in (msg_in_120), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u121 (.align_out (msg_out_121), .align_target_in (msg_in_121), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u122 (.align_out (msg_out_122), .align_target_in (msg_in_122), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u123 (.align_out (msg_out_123), .align_target_in (msg_in_123), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u124 (.align_out (msg_out_124), .align_target_in (msg_in_124), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u125 (.align_out (msg_out_125), .align_target_in (msg_in_125), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u126 (.align_out (msg_out_126), .align_target_in (msg_in_126), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u127 (.align_out (msg_out_127), .align_target_in (msg_in_127), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u128 (.align_out (msg_out_128), .align_target_in (msg_in_128), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u129 (.align_out (msg_out_129), .align_target_in (msg_in_129), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u130 (.align_out (msg_out_130), .align_target_in (msg_in_130), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u131 (.align_out (msg_out_131), .align_target_in (msg_in_131), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u132 (.align_out (msg_out_132), .align_target_in (msg_in_132), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u133 (.align_out (msg_out_133), .align_target_in (msg_in_133), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u134 (.align_out (msg_out_134), .align_target_in (msg_in_134), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u135 (.align_out (msg_out_135), .align_target_in (msg_in_135), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u136 (.align_out (msg_out_136), .align_target_in (msg_in_136), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u137 (.align_out (msg_out_137), .align_target_in (msg_in_137), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u138 (.align_out (msg_out_138), .align_target_in (msg_in_138), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u139 (.align_out (msg_out_139), .align_target_in (msg_in_139), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u140 (.align_out (msg_out_140), .align_target_in (msg_in_140), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u141 (.align_out (msg_out_141), .align_target_in (msg_in_141), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u142 (.align_out (msg_out_142), .align_target_in (msg_in_142), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u143 (.align_out (msg_out_143), .align_target_in (msg_in_143), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u144 (.align_out (msg_out_144), .align_target_in (msg_in_144), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u145 (.align_out (msg_out_145), .align_target_in (msg_in_145), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u146 (.align_out (msg_out_146), .align_target_in (msg_in_146), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u147 (.align_out (msg_out_147), .align_target_in (msg_in_147), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u148 (.align_out (msg_out_148), .align_target_in (msg_in_148), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u149 (.align_out (msg_out_149), .align_target_in (msg_in_149), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u150 (.align_out (msg_out_150), .align_target_in (msg_in_150), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u151 (.align_out (msg_out_151), .align_target_in (msg_in_151), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u152 (.align_out (msg_out_152), .align_target_in (msg_in_152), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u153 (.align_out (msg_out_153), .align_target_in (msg_in_153), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u154 (.align_out (msg_out_154), .align_target_in (msg_in_154), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u155 (.align_out (msg_out_155), .align_target_in (msg_in_155), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u156 (.align_out (msg_out_156), .align_target_in (msg_in_156), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u157 (.align_out (msg_out_157), .align_target_in (msg_in_157), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u158 (.align_out (msg_out_158), .align_target_in (msg_in_158), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u159 (.align_out (msg_out_159), .align_target_in (msg_in_159), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u160 (.align_out (msg_out_160), .align_target_in (msg_in_160), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u161 (.align_out (msg_out_161), .align_target_in (msg_in_161), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u162 (.align_out (msg_out_162), .align_target_in (msg_in_162), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u163 (.align_out (msg_out_163), .align_target_in (msg_in_163), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u164 (.align_out (msg_out_164), .align_target_in (msg_in_164), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u165 (.align_out (msg_out_165), .align_target_in (msg_in_165), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u166 (.align_out (msg_out_166), .align_target_in (msg_in_166), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u167 (.align_out (msg_out_167), .align_target_in (msg_in_167), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u168 (.align_out (msg_out_168), .align_target_in (msg_in_168), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u169 (.align_out (msg_out_169), .align_target_in (msg_in_169), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u170 (.align_out (msg_out_170), .align_target_in (msg_in_170), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u171 (.align_out (msg_out_171), .align_target_in (msg_in_171), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u172 (.align_out (msg_out_172), .align_target_in (msg_in_172), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u173 (.align_out (msg_out_173), .align_target_in (msg_in_173), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u174 (.align_out (msg_out_174), .align_target_in (msg_in_174), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u175 (.align_out (msg_out_175), .align_target_in (msg_in_175), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u176 (.align_out (msg_out_176), .align_target_in (msg_in_176), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u177 (.align_out (msg_out_177), .align_target_in (msg_in_177), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u178 (.align_out (msg_out_178), .align_target_in (msg_in_178), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u179 (.align_out (msg_out_179), .align_target_in (msg_in_179), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u180 (.align_out (msg_out_180), .align_target_in (msg_in_180), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u181 (.align_out (msg_out_181), .align_target_in (msg_in_181), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u182 (.align_out (msg_out_182), .align_target_in (msg_in_182), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u183 (.align_out (msg_out_183), .align_target_in (msg_in_183), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u184 (.align_out (msg_out_184), .align_target_in (msg_in_184), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u185 (.align_out (msg_out_185), .align_target_in (msg_in_185), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u186 (.align_out (msg_out_186), .align_target_in (msg_in_186), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u187 (.align_out (msg_out_187), .align_target_in (msg_in_187), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u188 (.align_out (msg_out_188), .align_target_in (msg_in_188), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u189 (.align_out (msg_out_189), .align_target_in (msg_in_189), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u190 (.align_out (msg_out_190), .align_target_in (msg_in_190), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u191 (.align_out (msg_out_191), .align_target_in (msg_in_191), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u192 (.align_out (msg_out_192), .align_target_in (msg_in_192), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u193 (.align_out (msg_out_193), .align_target_in (msg_in_193), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u194 (.align_out (msg_out_194), .align_target_in (msg_in_194), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u195 (.align_out (msg_out_195), .align_target_in (msg_in_195), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u196 (.align_out (msg_out_196), .align_target_in (msg_in_196), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u197 (.align_out (msg_out_197), .align_target_in (msg_in_197), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u198 (.align_out (msg_out_198), .align_target_in (msg_in_198), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u199 (.align_out (msg_out_199), .align_target_in (msg_in_199), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u200 (.align_out (msg_out_200), .align_target_in (msg_in_200), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u201 (.align_out (msg_out_201), .align_target_in (msg_in_201), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u202 (.align_out (msg_out_202), .align_target_in (msg_in_202), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u203 (.align_out (msg_out_203), .align_target_in (msg_in_203), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u204 (.align_out (msg_out_204), .align_target_in (msg_in_204), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u205 (.align_out (msg_out_205), .align_target_in (msg_in_205), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u206 (.align_out (msg_out_206), .align_target_in (msg_in_206), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u207 (.align_out (msg_out_207), .align_target_in (msg_in_207), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u208 (.align_out (msg_out_208), .align_target_in (msg_in_208), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u209 (.align_out (msg_out_209), .align_target_in (msg_in_209), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u210 (.align_out (msg_out_210), .align_target_in (msg_in_210), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u211 (.align_out (msg_out_211), .align_target_in (msg_in_211), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u212 (.align_out (msg_out_212), .align_target_in (msg_in_212), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u213 (.align_out (msg_out_213), .align_target_in (msg_in_213), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u214 (.align_out (msg_out_214), .align_target_in (msg_in_214), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u215 (.align_out (msg_out_215), .align_target_in (msg_in_215), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u216 (.align_out (msg_out_216), .align_target_in (msg_in_216), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u217 (.align_out (msg_out_217), .align_target_in (msg_in_217), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u218 (.align_out (msg_out_218), .align_target_in (msg_in_218), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u219 (.align_out (msg_out_219), .align_target_in (msg_in_219), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u220 (.align_out (msg_out_220), .align_target_in (msg_in_220), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u221 (.align_out (msg_out_221), .align_target_in (msg_in_221), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u222 (.align_out (msg_out_222), .align_target_in (msg_in_222), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u223 (.align_out (msg_out_223), .align_target_in (msg_in_223), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u224 (.align_out (msg_out_224), .align_target_in (msg_in_224), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u225 (.align_out (msg_out_225), .align_target_in (msg_in_225), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u226 (.align_out (msg_out_226), .align_target_in (msg_in_226), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u227 (.align_out (msg_out_227), .align_target_in (msg_in_227), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u228 (.align_out (msg_out_228), .align_target_in (msg_in_228), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u229 (.align_out (msg_out_229), .align_target_in (msg_in_229), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u230 (.align_out (msg_out_230), .align_target_in (msg_in_230), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u231 (.align_out (msg_out_231), .align_target_in (msg_in_231), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u232 (.align_out (msg_out_232), .align_target_in (msg_in_232), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u233 (.align_out (msg_out_233), .align_target_in (msg_in_233), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u234 (.align_out (msg_out_234), .align_target_in (msg_in_234), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u235 (.align_out (msg_out_235), .align_target_in (msg_in_235), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u236 (.align_out (msg_out_236), .align_target_in (msg_in_236), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u237 (.align_out (msg_out_237), .align_target_in (msg_in_237), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u238 (.align_out (msg_out_238), .align_target_in (msg_in_238), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u239 (.align_out (msg_out_239), .align_target_in (msg_in_239), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u240 (.align_out (msg_out_240), .align_target_in (msg_in_240), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u241 (.align_out (msg_out_241), .align_target_in (msg_in_241), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u242 (.align_out (msg_out_242), .align_target_in (msg_in_242), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u243 (.align_out (msg_out_243), .align_target_in (msg_in_243), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u244 (.align_out (msg_out_244), .align_target_in (msg_in_244), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u245 (.align_out (msg_out_245), .align_target_in (msg_in_245), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u246 (.align_out (msg_out_246), .align_target_in (msg_in_246), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u247 (.align_out (msg_out_247), .align_target_in (msg_in_247), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u248 (.align_out (msg_out_248), .align_target_in (msg_in_248), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u249 (.align_out (msg_out_249), .align_target_in (msg_in_249), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u250 (.align_out (msg_out_250), .align_target_in (msg_in_250), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u251 (.align_out (msg_out_251), .align_target_in (msg_in_251), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u252 (.align_out (msg_out_252), .align_target_in (msg_in_252), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u253 (.align_out (msg_out_253), .align_target_in (msg_in_253), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
circular_page_align_depth_1 #(.QUAN_SIZE (QUAN_SIZE)) page_align_u254 (.align_out (msg_out_254), .align_target_in (msg_in_254), .first_row_chunk(first_row_chunk), .sys_clk(sys_clk), .rstn(rstn));
/////////////////////////////////////////////////////////////////////////////////////////////
endmodule
`endif